* File created on: 2025-05-09 14:30:08
* From this circuit description: ../../examples/INV_string_11_CC_RBUS_SBUS.json
* "spice" description for "MOSbius_v2_tb", "PK_set_SWMATRIX", "spice" 


simulator lang=spice

.SUBCKT PK_set_SWMATRIX PROBE<1> PROBE<2> PROBE<3> PROBE<4> PROBE<5> PROBE<6>
+  PROBE<7> PROBE<8> PROBE<9> PROBE<10> PROBE<11> PROBE<12> PROBE<13> PROBE<14>
+  PROBE<15> PROBE<16> PROBE<17> PROBE<18> PROBE<19> PROBE<20> PROBE<21>
+  PROBE<22> PROBE<23> PROBE<24> PROBE<25> PROBE<26> PROBE<27> PROBE<28>
+  PROBE<29> PROBE<30> PROBE<31> PROBE<32> PROBE<33> PROBE<34> PROBE<35>
+  PROBE<36> PROBE<37> PROBE<38> PROBE<39> PROBE<40> PROBE<41> PROBE<42>
+  PROBE<43> PROBE<44> PROBE<45> PROBE<46> PROBE<47> PROBE<48> PROBE<49>
+  PROBE<50> PROBE<51> PROBE<52> PROBE<53> PROBE<54> PROBE<55> PROBE<56>
+  PROBE<57> PROBE<58> PROBE<59> PROBE<60> PROBE<61> PROBE<62> PROBE<63>
+  PROBE<64> PROBE<65> PROBE<66> PROBE<67> PROBE<68> PROBE<69> PROBE<70>
+  PROBE<71> PROBE<72> PROBE<73> PROBE<74> PROBE<75> PROBE<76> PROBE<77>
+  PROBE<78> PROBE<79> PROBE<80> PROBE<81> PROBE<82> PROBE<83> PROBE<84>
+  PROBE<85> PROBE<86> PROBE<87> PROBE<88> PROBE<89> PROBE<90> PROBE<91>
+  PROBE<92> PROBE<93> PROBE<94> PROBE<95> PROBE<96> PROBE<97> PROBE<98>
+  PROBE<99> PROBE<100> PROBE<101> PROBE<102> PROBE<103> PROBE<104> PROBE<105>
+  PROBE<106> PROBE<107> PROBE<108> PROBE<109> PROBE<110> PROBE<111> PROBE<112>
+  PROBE<113> PROBE<114> PROBE<115> PROBE<116> PROBE<117> PROBE<118> PROBE<119>
+  PROBE<120> PROBE<121> PROBE<122> PROBE<123> PROBE<124> PROBE<125> PROBE<126>
+  PROBE<127> PROBE<128> PROBE<129> PROBE<130> PROBE<131> PROBE<132> PROBE<133>
+  PROBE<134> PROBE<135> PROBE<136> PROBE<137> PROBE<138> PROBE<139> PROBE<140>
+  PROBE<141> PROBE<142> PROBE<143> PROBE<144> PROBE<145> PROBE<146> PROBE<147>
+  PROBE<148> PROBE<149> PROBE<150> PROBE<151> PROBE<152> PROBE<153> PROBE<154>
+  PROBE<155> PROBE<156> PROBE<157> PROBE<158> PROBE<159> PROBE<160> PROBE<161>
+  PROBE<162> PROBE<163> PROBE<164> PROBE<165> PROBE<166> PROBE<167> PROBE<168>
+  PROBE<169> PROBE<170> PROBE<171> PROBE<172> PROBE<173> PROBE<174> PROBE<175>
+  PROBE<176> PROBE<177> PROBE<178> PROBE<179> PROBE<180> PROBE<181> PROBE<182>
+  PROBE<183> PROBE<184> PROBE<185> PROBE<186> PROBE<187> PROBE<188> PROBE<189>
+  PROBE<190> PROBE<191> PROBE<192> PROBE<193> PROBE<194> PROBE<195> PROBE<196>
+  PROBE<197> PROBE<198> PROBE<199> PROBE<200> PROBE<201> PROBE<202> PROBE<203>
+  PROBE<204> PROBE<205> PROBE<206> PROBE<207> PROBE<208> PROBE<209> PROBE<210>
+  PROBE<211> PROBE<212> PROBE<213> PROBE<214> PROBE<215> PROBE<216> PROBE<217>
+  PROBE<218> PROBE<219> PROBE<220> PROBE<221> PROBE<222> PROBE<223> PROBE<224>
+  PROBE<225> PROBE<226> PROBE<227> PROBE<228> PROBE<229> PROBE<230> PROBE<231>
+  PROBE<232> PROBE<233> PROBE<234> PROBE<235> PROBE<236> PROBE<237> PROBE<238>
+  PROBE<239> PROBE<240> PROBE<241> PROBE<242> PROBE<243> PROBE<244> PROBE<245>
+  PROBE<246> PROBE<247> PROBE<248> PROBE<249> PROBE<250> PROBE<251> PROBE<252>
+  PROBE<253> PROBE<254> PROBE<255> PROBE<256> PROBE<257> PROBE<258> PROBE<259>
+  PROBE<260> PROBE<261> PROBE<262> PROBE<263> PROBE<264> PROBE<265> PROBE<266>
+  PROBE<267> PROBE<268> PROBE<269> PROBE<270> PROBE<271> PROBE<272> PROBE<273>
+  PROBE<274> PROBE<275> PROBE<276> PROBE<277> PROBE<278> PROBE<279> PROBE<280>
+  PROBE<281> PROBE<282> PROBE<283> PROBE<284> PROBE<285> PROBE<286> PROBE<287>
+  PROBE<288> PROBE<289> PROBE<290> PROBE<291> PROBE<292> PROBE<293> PROBE<294>
+  PROBE<295> PROBE<296> PROBE<297> PROBE<298> PROBE<299> PROBE<300> PROBE<301>
+  PROBE<302> PROBE<303> PROBE<304> PROBE<305> PROBE<306> PROBE<307> PROBE<308>
+  PROBE<309> PROBE<310> PROBE<311> PROBE<312> PROBE<313> PROBE<314> PROBE<315>
+  PROBE<316> PROBE<317> PROBE<318> PROBE<319> PROBE<320> PROBE<321> PROBE<322>
+  PROBE<323> PROBE<324> PROBE<325> PROBE<326> PROBE<327> PROBE<328> PROBE<329>
+  PROBE<330> PROBE<331> PROBE<332> PROBE<333> PROBE<334> PROBE<335> PROBE<336>
+  PROBE<337> PROBE<338> PROBE<339> PROBE<340> PROBE<341> PROBE<342> PROBE<343>
+  PROBE<344> PROBE<345> PROBE<346> PROBE<347> PROBE<348> PROBE<349> PROBE<350>
+  PROBE<351> PROBE<352> PROBE<353> PROBE<354> PROBE<355> PROBE<356> PROBE<357>
+  PROBE<358> PROBE<359> PROBE<360> PROBE<361> PROBE<362> PROBE<363> PROBE<364>
+  PROBE<365> PROBE<366> PROBE<367> PROBE<368> PROBE<369> PROBE<370> PROBE<371>
+  PROBE<372> PROBE<373> PROBE<374> PROBE<375> PROBE<376> PROBE<377> PROBE<378>
+  PROBE<379> PROBE<380> PROBE<381> PROBE<382> PROBE<383> PROBE<384> PROBE<385>
+  PROBE<386> PROBE<387> PROBE<388> PROBE<389> PROBE<390> PROBE<391> PROBE<392>
+  PROBE<393> PROBE<394> PROBE<395> PROBE<396> PROBE<397> PROBE<398> PROBE<399>
+  PROBE<400> PROBE<401> PROBE<402> PROBE<403> PROBE<404> PROBE<405> PROBE<406>
+  PROBE<407> PROBE<408> PROBE<409> PROBE<410> PROBE<411> PROBE<412> PROBE<413>
+  PROBE<414> PROBE<415> PROBE<416> PROBE<417> PROBE<418> PROBE<419> PROBE<420>
+  PROBE<421> PROBE<422> PROBE<423> PROBE<424> PROBE<425> PROBE<426> PROBE<427>
+  PROBE<428> PROBE<429> PROBE<430> PROBE<431> PROBE<432> PROBE<433> PROBE<434>
+  PROBE<435> PROBE<436> PROBE<437> PROBE<438> PROBE<439> PROBE<440> PROBE<441>
+  PROBE<442> PROBE<443> PROBE<444> PROBE<445> PROBE<446> PROBE<447> PROBE<448>
+  PROBE<449> PROBE<450> PROBE<451> PROBE<452> PROBE<453> PROBE<454> PROBE<455>
+  PROBE<456> PROBE<457> PROBE<458> PROBE<459> PROBE<460> PROBE<461> PROBE<462>
+  PROBE<463> PROBE<464> PROBE<465> PROBE<466> PROBE<467> PROBE<468> PROBE<469>
+  PROBE<470> PROBE<471> PROBE<472> PROBE<473> PROBE<474> PROBE<475> PROBE<476>
+  PROBE<477> PROBE<478> PROBE<479> PROBE<480> PROBE<481> PROBE<482> PROBE<483>
+  PROBE<484> PROBE<485> PROBE<486> PROBE<487> PROBE<488> PROBE<489> PROBE<490>
+  PROBE<491> PROBE<492> PROBE<493> PROBE<494> PROBE<495> PROBE<496> PROBE<497>
+  PROBE<498> PROBE<499> PROBE<500> PROBE<501> PROBE<502> PROBE<503> PROBE<504>
+  PROBE<505> PROBE<506> PROBE<507> PROBE<508> PROBE<509> PROBE<510> PROBE<511>
+  PROBE<512> PROBE<513> PROBE<514> PROBE<515> PROBE<516> PROBE<517> PROBE<518>
+  PROBE<519> PROBE<520> PROBE<521> PROBE<522> PROBE<523> PROBE<524> PROBE<525>
+  PROBE<526> PROBE<527> PROBE<528> PROBE<529> PROBE<530> PROBE<531> PROBE<532>
+  PROBE<533> PROBE<534> PROBE<535> PROBE<536> PROBE<537> PROBE<538> PROBE<539>
+  PROBE<540> PROBE<541> PROBE<542> PROBE<543> PROBE<544> PROBE<545> PROBE<546>
+  PROBE<547> PROBE<548> PROBE<549> PROBE<550> PROBE<551> PROBE<552> PROBE<553>
+  PROBE<554> PROBE<555> PROBE<556> PROBE<557> PROBE<558> PROBE<559> PROBE<560>
+  PROBE<561> PROBE<562> PROBE<563> PROBE<564> PROBE<565> PROBE<566> PROBE<567>
+  PROBE<568> PROBE<569> PROBE<570> PROBE<571> PROBE<572> PROBE<573> PROBE<574>
+  PROBE<575> PROBE<576> PROBE<577> PROBE<578> PROBE<579> PROBE<580> PROBE<581>
+  PROBE<582> PROBE<583> PROBE<584> PROBE<585> PROBE<586> PROBE<587> PROBE<588>
+  PROBE<589> PROBE<590> PROBE<591> PROBE<592> PROBE<593> PROBE<594> PROBE<595>
+  PROBE<596> PROBE<597> PROBE<598> PROBE<599> PROBE<600> PROBE<601> PROBE<602>
+  PROBE<603> PROBE<604> PROBE<605> PROBE<606> PROBE<607> PROBE<608> PROBE<609>
+  PROBE<610> PROBE<611> PROBE<612> PROBE<613> PROBE<614> PROBE<615> PROBE<616>
+  PROBE<617> PROBE<618> PROBE<619> PROBE<620> PROBE<621> PROBE<622> PROBE<623>
+  PROBE<624> PROBE<625> PROBE<626> PROBE<627> PROBE<628> PROBE<629> PROBE<630>
+  PROBE<631> PROBE<632> PROBE<633> PROBE<634> PROBE<635> PROBE<636> PROBE<637>
+  PROBE<638> PROBE<639> PROBE<640> PROBE<641> PROBE<642> PROBE<643> PROBE<644>
+  PROBE<645> PROBE<646> PROBE<647> PROBE<648> PROBE<649> PROBE<650> PROBE<651>
+  PROBE<652> PROBE<653> PROBE<654> PROBE<655> PROBE<656> PROBE<657> PROBE<658>
+  PROBE<659> PROBE<660> PROBE<661> PROBE<662> PROBE<663> PROBE<664> PROBE<665>
+  PROBE<666> PROBE<667> PROBE<668> PROBE<669> PROBE<670> PROBE<671> PROBE<672>
+  PROBE<673> PROBE<674> PROBE<675> PROBE<676> PROBE<677> PROBE<678> PROBE<679>
+  PROBE<680> PROBE<681> PROBE<682> PROBE<683> PROBE<684> PROBE<685> PROBE<686>
+  PROBE<687> PROBE<688> PROBE<689> PROBE<690> PROBE<691> PROBE<692> PROBE<693>
+  PROBE<694> PROBE<695> PROBE<696> PROBE<697> PROBE<698> PROBE<699> PROBE<700>
+  PROBE<701> PROBE<702> PROBE<703> PROBE<704> PROBE<705> PROBE<706> PROBE<707>
+  PROBE<708> PROBE<709> PROBE<710> PROBE<711> PROBE<712> PROBE<713> PROBE<714>
+  PROBE<715> PROBE<716> PROBE<717> PROBE<718> PROBE<719> PROBE<720> PROBE<721>
+  PROBE<722> PROBE<723> PROBE<724> PROBE<725> PROBE<726> PROBE<727> PROBE<728>
+  PROBE<729> PROBE<730> PROBE<731> PROBE<732> PROBE<733> PROBE<734> PROBE<735>
+  PROBE<736> PROBE<737> PROBE<738> PROBE<739> PROBE<740> PROBE<741> PROBE<742>
+  PROBE<743> PROBE<744> PROBE<745> PROBE<746> PROBE<747> PROBE<748> PROBE<749>
+  PROBE<750> PROBE<751> PROBE<752> PROBE<753> PROBE<754> PROBE<755> PROBE<756>
+  PROBE<757> PROBE<758> PROBE<759> PROBE<760> PROBE<761> PROBE<762> PROBE<763>
+  PROBE<764> PROBE<765> PROBE<766> PROBE<767> PROBE<768> PROBE<769> PROBE<770>
+  PROBE<771> PROBE<772> PROBE<773> PROBE<774> PROBE<775> PROBE<776> PROBE<777>
+  PROBE<778> PROBE<779> PROBE<780> PROBE<781> PROBE<782> PROBE<783> PROBE<784>
+  PROBE<785> PROBE<786> PROBE<787> PROBE<788> PROBE<789> PROBE<790> PROBE<791>
+  PROBE<792> PROBE<793> PROBE<794> PROBE<795> PROBE<796> PROBE<797> PROBE<798>
+  PROBE<799> PROBE<800> PROBE<801> PROBE<802> PROBE<803> PROBE<804> PROBE<805>
+  PROBE<806> PROBE<807> PROBE<808> PROBE<809> PROBE<810> PROBE<811> PROBE<812>
+  PROBE<813> PROBE<814> PROBE<815> PROBE<816> PROBE<817> PROBE<818> PROBE<819>
+  PROBE<820> PROBE<821> PROBE<822> PROBE<823> PROBE<824> PROBE<825> PROBE<826>
+  PROBE<827> PROBE<828> PROBE<829> PROBE<830> PROBE<831> PROBE<832> PROBE<833>
+  PROBE<834> PROBE<835> PROBE<836> PROBE<837> PROBE<838> PROBE<839> PROBE<840>
+  PROBE<841> PROBE<842> PROBE<843> PROBE<844> PROBE<845> PROBE<846> PROBE<847>
+  PROBE<848> PROBE<849> PROBE<850> PROBE<851> PROBE<852> PROBE<853> PROBE<854>
+  PROBE<855> PROBE<856> PROBE<857> PROBE<858> PROBE<859> PROBE<860> PROBE<861>
+  PROBE<862> PROBE<863> PROBE<864> PROBE<865> PROBE<866> PROBE<867> PROBE<868>
+  PROBE<869> PROBE<870> PROBE<871> PROBE<872> PROBE<873> PROBE<874> PROBE<875>
+  PROBE<876> PROBE<877> PROBE<878> PROBE<879> PROBE<880> PROBE<881> PROBE<882>
+  PROBE<883> PROBE<884> PROBE<885> PROBE<886> PROBE<887> PROBE<888> PROBE<889>
+  PROBE<890> PROBE<891> PROBE<892> PROBE<893> PROBE<894> PROBE<895> PROBE<896>
+  PROBE<897> PROBE<898> PROBE<899> PROBE<900> PROBE<901> PROBE<902> PROBE<903>
+  PROBE<904> PROBE<905> PROBE<906> PROBE<907> PROBE<908> PROBE<909> PROBE<910>
+  PROBE<911> PROBE<912> PROBE<913> PROBE<914> PROBE<915> PROBE<916> PROBE<917>
+  PROBE<918> PROBE<919> PROBE<920> PROBE<921> PROBE<922> PROBE<923> PROBE<924>
+  PROBE<925> PROBE<926> PROBE<927> PROBE<928> PROBE<929> PROBE<930> PROBE<931>
+  PROBE<932> PROBE<933> PROBE<934> PROBE<935> PROBE<936> PROBE<937> PROBE<938>
+  PROBE<939> PROBE<940> PROBE<941> PROBE<942> PROBE<943> PROBE<944> PROBE<945>
+  PROBE<946> PROBE<947> PROBE<948> PROBE<949> PROBE<950> PROBE<951> PROBE<952>
+  PROBE<953> PROBE<954> PROBE<955> PROBE<956> PROBE<957> PROBE<958> PROBE<959>
+  PROBE<960> PROBE<961> PROBE<962> PROBE<963> PROBE<964> PROBE<965> PROBE<966>
+  PROBE<967> PROBE<968> PROBE<969> PROBE<970> PROBE<971> PROBE<972> PROBE<973>
+  PROBE<974> PROBE<975> PROBE<976> PROBE<977> PROBE<978> PROBE<979> PROBE<980>
+  PROBE<981> PROBE<982> PROBE<983> PROBE<984> PROBE<985> PROBE<986> PROBE<987>
+  PROBE<988> PROBE<989> PROBE<990> PROBE<991> PROBE<992> PROBE<993> PROBE<994>
+  PROBE<995> PROBE<996> PROBE<997> PROBE<998> PROBE<999> PROBE<1000> PROBE<1001>
+  PROBE<1002> PROBE<1003> PROBE<1004> PROBE<1005> PROBE<1006> PROBE<1007>
+  PROBE<1008> PROBE<1009> PROBE<1010> PROBE<1011> PROBE<1012> PROBE<1013>
+  PROBE<1014> PROBE<1015> PROBE<1016> PROBE<1017> PROBE<1018> PROBE<1019>
+  PROBE<1020> PROBE<1021> PROBE<1022> PROBE<1023> PROBE<1024> PROBE<1025>
+  PROBE<1026> PROBE<1027> PROBE<1028> PROBE<1029> PROBE<1030> PROBE<1031>
+  PROBE<1032> PROBE<1033> PROBE<1034> PROBE<1035> PROBE<1036> PROBE<1037>
+  PROBE<1038> PROBE<1039> PROBE<1040> PROBE<1041> PROBE<1042> PROBE<1043>
+  PROBE<1044> PROBE<1045> PROBE<1046> PROBE<1047> PROBE<1048> PROBE<1049>
+  PROBE<1050> PROBE<1051> PROBE<1052> PROBE<1053> PROBE<1054> PROBE<1055>
+  PROBE<1056> PROBE<1057> PROBE<1058> PROBE<1059> PROBE<1060> PROBE<1061>
+  PROBE<1062> PROBE<1063> PROBE<1064> PROBE<1065> PROBE<1066> PROBE<1067>
+  PROBE<1068> PROBE<1069> PROBE<1070> PROBE<1071> PROBE<1072> PROBE<1073>
+  PROBE<1074> PROBE<1075> PROBE<1076> PROBE<1077> PROBE<1078> PROBE<1079>
+  PROBE<1080> PROBE<1081> PROBE<1082> PROBE<1083> PROBE<1084> PROBE<1085>
+  PROBE<1086> PROBE<1087> PROBE<1088> PROBE<1089> PROBE<1090> PROBE<1091>
+  PROBE<1092> PROBE<1093> PROBE<1094> PROBE<1095> PROBE<1096> PROBE<1097>
+  PROBE<1098> PROBE<1099> PROBE<1100> PROBE<1101> PROBE<1102> PROBE<1103>
+  PROBE<1104> PROBE<1105> PROBE<1106> PROBE<1107> PROBE<1108> PROBE<1109>
+  PROBE<1110> PROBE<1111> PROBE<1112> PROBE<1113> PROBE<1114> PROBE<1115>
+  PROBE<1116> PROBE<1117> PROBE<1118> PROBE<1119> PROBE<1120> PROBE<1121>
+  PROBE<1122> PROBE<1123> PROBE<1124> PROBE<1125> PROBE<1126> PROBE<1127>
+  PROBE<1128> PROBE<1129> PROBE<1130> PROBE<1131> PROBE<1132> PROBE<1133>
+  PROBE<1134> PROBE<1135> PROBE<1136> PROBE<1137> PROBE<1138> PROBE<1139>
+  PROBE<1140> PROBE<1141> PROBE<1142> PROBE<1143> PROBE<1144> PROBE<1145>
+  PROBE<1146> PROBE<1147> PROBE<1148> PROBE<1149> PROBE<1150> PROBE<1151>
+  PROBE<1152> PROBE<1153> PROBE<1154> PROBE<1155> PROBE<1156> PROBE<1157>
+  PROBE<1158> PROBE<1159> PROBE<1160> PROBE<1161> PROBE<1162> PROBE<1163>
+  PROBE<1164> PROBE<1165> PROBE<1166> PROBE<1167> PROBE<1168> PROBE<1169>
+  PROBE<1170> PROBE<1171> PROBE<1172> PROBE<1173> PROBE<1174> PROBE<1175>
+  PROBE<1176> PROBE<1177> PROBE<1178> PROBE<1179> PROBE<1180> PROBE<1181>
+  PROBE<1182> PROBE<1183> PROBE<1184> PROBE<1185> PROBE<1186> PROBE<1187>
+  PROBE<1188> PROBE<1189> PROBE<1190> PROBE<1191> PROBE<1192> PROBE<1193>
+  PROBE<1194> PROBE<1195> PROBE<1196> PROBE<1197> PROBE<1198> PROBE<1199>
+  PROBE<1200> PROBE<1201> PROBE<1202> PROBE<1203> PROBE<1204> PROBE<1205>
+  PROBE<1206> PROBE<1207> PROBE<1208> PROBE<1209> PROBE<1210> PROBE<1211>
+  PROBE<1212> PROBE<1213> PROBE<1214> PROBE<1215> PROBE<1216> PROBE<1217>
+  PROBE<1218> PROBE<1219> PROBE<1220> PROBE<1221> PROBE<1222> PROBE<1223>
+  PROBE<1224> PROBE<1225> PROBE<1226> PROBE<1227> PROBE<1228> PROBE<1229>
+  PROBE<1230> PROBE<1231> PROBE<1232> PROBE<1233> PROBE<1234> PROBE<1235>
+  PROBE<1236> PROBE<1237> PROBE<1238> PROBE<1239> PROBE<1240> PROBE<1241>
+  PROBE<1242> PROBE<1243> PROBE<1244> PROBE<1245> PROBE<1246> PROBE<1247>
+  PROBE<1248> PROBE<1249> PROBE<1250> PROBE<1251> PROBE<1252> PROBE<1253>
+  PROBE<1254> PROBE<1255> PROBE<1256> PROBE<1257> PROBE<1258> PROBE<1259>
+  PROBE<1260> PROBE<1261> PROBE<1262> PROBE<1263> PROBE<1264> PROBE<1265>
+  PROBE<1266> PROBE<1267> PROBE<1268> PROBE<1269> PROBE<1270> PROBE<1271>
+  PROBE<1272> PROBE<1273> PROBE<1274> PROBE<1275> PROBE<1276> PROBE<1277>
+  PROBE<1278> PROBE<1279> PROBE<1280> PROBE<1281> PROBE<1282> PROBE<1283>
+  PROBE<1284> PROBE<1285> PROBE<1286> PROBE<1287> PROBE<1288> PROBE<1289>
+  PROBE<1290> PROBE<1291> PROBE<1292> PROBE<1293> PROBE<1294> PROBE<1295>
+  PROBE<1296> PROBE<1297> PROBE<1298> PROBE<1299> PROBE<1300> PROBE<1301>
+  PROBE<1302> PROBE<1303> PROBE<1304> PROBE<1305> PROBE<1306> PROBE<1307>
+  PROBE<1308> PROBE<1309> PROBE<1310> PROBE<1311> PROBE<1312> PROBE<1313>
+  PROBE<1314> PROBE<1315> PROBE<1316> PROBE<1317> PROBE<1318> PROBE<1319>
+  PROBE<1320> PROBE<1321> PROBE<1322> PROBE<1323> PROBE<1324> PROBE<1325>
+  PROBE<1326> PROBE<1327> PROBE<1328> PROBE<1329> PROBE<1330> PROBE<1331>
+  PROBE<1332> PROBE<1333> PROBE<1334> PROBE<1335> PROBE<1336> PROBE<1337>
+  PROBE<1338> PROBE<1339> PROBE<1340> PROBE<1341> PROBE<1342> PROBE<1343>
+  PROBE<1344> PROBE<1345> PROBE<1346> PROBE<1347> PROBE<1348> PROBE<1349>
+  PROBE<1350> PROBE<1351> PROBE<1352> PROBE<1353> PROBE<1354> PROBE<1355>
+  PROBE<1356> PROBE<1357> PROBE<1358> PROBE<1359> PROBE<1360> PROBE<1361>
+  PROBE<1362> PROBE<1363> PROBE<1364> PROBE<1365> PROBE<1366> PROBE<1367>
+  PROBE<1368> PROBE<1369> PROBE<1370> PROBE<1371> PROBE<1372> PROBE<1373>
+  PROBE<1374> PROBE<1375> PROBE<1376> PROBE<1377> PROBE<1378> PROBE<1379>
+  PROBE<1380> PROBE<1381> PROBE<1382> PROBE<1383> PROBE<1384> PROBE<1385>
+  PROBE<1386> PROBE<1387> PROBE<1388> PROBE<1389> PROBE<1390> PROBE<1391>
+  PROBE<1392> PROBE<1393> PROBE<1394> PROBE<1395> PROBE<1396> PROBE<1397>
+  PROBE<1398> PROBE<1399> PROBE<1400> PROBE<1401> PROBE<1402> PROBE<1403>
+  PROBE<1404> PROBE<1405> PROBE<1406> PROBE<1407> PROBE<1408> PROBE<1409>
+  PROBE<1410> PROBE<1411> PROBE<1412> PROBE<1413> PROBE<1414> PROBE<1415>
+  PROBE<1416> PROBE<1417> PROBE<1418> PROBE<1419> PROBE<1420> PROBE<1421>
+  PROBE<1422> PROBE<1423> PROBE<1424> PROBE<1425> PROBE<1426> PROBE<1427>
+  PROBE<1428> PROBE<1429> PROBE<1430> PROBE<1431> PROBE<1432> PROBE<1433>
+  PROBE<1434> PROBE<1435> PROBE<1436> PROBE<1437> PROBE<1438> PROBE<1439>
+  PROBE<1440> PROBE<1441> PROBE<1442> PROBE<1443> PROBE<1444> PROBE<1445>
+  PROBE<1446> PROBE<1447> PROBE<1448> PROBE<1449> PROBE<1450> PROBE<1451>
+  PROBE<1452> PROBE<1453> PROBE<1454> PROBE<1455> PROBE<1456> PROBE<1457>
+  PROBE<1458> PROBE<1459> PROBE<1460> PROBE<1461> PROBE<1462> PROBE<1463>
+  PROBE<1464> PROBE<1465> PROBE<1466> PROBE<1467> PROBE<1468> PROBE<1469>
+  PROBE<1470> PROBE<1471> PROBE<1472> PROBE<1473> PROBE<1474> PROBE<1475>
+  PROBE<1476> PROBE<1477> PROBE<1478> PROBE<1479> PROBE<1480> PROBE<1481>
+  PROBE<1482> PROBE<1483> PROBE<1484> PROBE<1485> PROBE<1486> PROBE<1487>
+  PROBE<1488> PROBE<1489> PROBE<1490> PROBE<1491> PROBE<1492> PROBE<1493>
+  PROBE<1494> PROBE<1495> PROBE<1496> PROBE<1497> PROBE<1498> PROBE<1499>
+  PROBE<1500> PROBE<1501> PROBE<1502> PROBE<1503> PROBE<1504> PROBE<1505>
+  PROBE<1506> PROBE<1507> PROBE<1508> PROBE<1509> PROBE<1510> PROBE<1511>
+  PROBE<1512> PROBE<1513> PROBE<1514> PROBE<1515> PROBE<1516> PROBE<1517>
+  PROBE<1518> PROBE<1519> PROBE<1520> PROBE<1521> PROBE<1522> PROBE<1523>
+  PROBE<1524> PROBE<1525> PROBE<1526> PROBE<1527> PROBE<1528> PROBE<1529>
+  PROBE<1530> PROBE<1531> PROBE<1532> PROBE<1533> PROBE<1534> PROBE<1535>
+  PROBE<1536> PROBE<1537> PROBE<1538> PROBE<1539> PROBE<1540> PROBE<1541>
+  PROBE<1542> PROBE<1543> PROBE<1544> PROBE<1545> PROBE<1546> PROBE<1547>
+  PROBE<1548> PROBE<1549> PROBE<1550> PROBE<1551> PROBE<1552> PROBE<1553>
+  PROBE<1554> PROBE<1555> PROBE<1556> PROBE<1557> PROBE<1558> PROBE<1559>
+  PROBE<1560> PROBE<1561> PROBE<1562> PROBE<1563> PROBE<1564> PROBE<1565>
+  PROBE<1566> PROBE<1567> PROBE<1568> PROBE<1569> PROBE<1570> PROBE<1571>
+  PROBE<1572> PROBE<1573> PROBE<1574> PROBE<1575> PROBE<1576> PROBE<1577>
+  PROBE<1578> PROBE<1579> PROBE<1580> PROBE<1581> PROBE<1582> PROBE<1583>
+  PROBE<1584> PROBE<1585> PROBE<1586> PROBE<1587> PROBE<1588> PROBE<1589>
+  PROBE<1590> PROBE<1591> PROBE<1592> PROBE<1593> PROBE<1594> PROBE<1595>
+  PROBE<1596> PROBE<1597> PROBE<1598> PROBE<1599> PROBE<1600> PROBE<1601>
+  PROBE<1602> PROBE<1603> PROBE<1604> PROBE<1605> PROBE<1606> PROBE<1607>
+  PROBE<1608> PROBE<1609> PROBE<1610> PROBE<1611> PROBE<1612> PROBE<1613>
+  PROBE<1614> PROBE<1615> PROBE<1616> PROBE<1617> PROBE<1618> PROBE<1619>
+  PROBE<1620> PROBE<1621> PROBE<1622> PROBE<1623> PROBE<1624> PROBE<1625>
+  PROBE<1626> PROBE<1627> PROBE<1628> PROBE<1629> PROBE<1630> PROBE<1631>
+  PROBE<1632> PROBE<1633> PROBE<1634> PROBE<1635> PROBE<1636> PROBE<1637>
+  PROBE<1638> PROBE<1639> PROBE<1640> PROBE<1641> PROBE<1642> PROBE<1643>
+  PROBE<1644> PROBE<1645> PROBE<1646> PROBE<1647> PROBE<1648> PROBE<1649>
+  PROBE<1650> PROBE<1651> PROBE<1652> PROBE<1653> PROBE<1654> PROBE<1655>
+  PROBE<1656> PROBE<1657> PROBE<1658> PROBE<1659> PROBE<1660> PROBE<1661>
+  PROBE<1662> PROBE<1663> PROBE<1664> PROBE<1665> PROBE<1666> PROBE<1667>
+  PROBE<1668> PROBE<1669> PROBE<1670> PROBE<1671> PROBE<1672> PROBE<1673>
+  PROBE<1674> PROBE<1675> PROBE<1676> PROBE<1677> PROBE<1678> PROBE<1679>
+  PROBE<1680> PROBE<1681> PROBE<1682> PROBE<1683> PROBE<1684> PROBE<1685>
+  PROBE<1686> PROBE<1687> PROBE<1688> PROBE<1689> PROBE<1690> PROBE<1691>
+  PROBE<1692> PROBE<1693> PROBE<1694> PROBE<1695> PROBE<1696> PROBE<1697>
+  PROBE<1698> PROBE<1699> PROBE<1700> PROBE<1701> PROBE<1702> PROBE<1703>
+  PROBE<1704> PROBE<1705> PROBE<1706> PROBE<1707> PROBE<1708> PROBE<1709>
+  PROBE<1710> PROBE<1711> PROBE<1712> PROBE<1713> PROBE<1714> PROBE<1715>
+  PROBE<1716> PROBE<1717> PROBE<1718> PROBE<1719> PROBE<1720> PROBE<1721>
+  PROBE<1722> PROBE<1723> PROBE<1724> PROBE<1725> PROBE<1726> PROBE<1727>
+  PROBE<1728> PROBE<1729> PROBE<1730> PROBE<1731> PROBE<1732> PROBE<1733>
+  PROBE<1734> PROBE<1735> PROBE<1736> PROBE<1737> PROBE<1738> PROBE<1739>
+  PROBE<1740> PROBE<1741> PROBE<1742> PROBE<1743> PROBE<1744> PROBE<1745>
+  PROBE<1746> PROBE<1747> PROBE<1748> PROBE<1749> PROBE<1750> PROBE<1751>
+  PROBE<1752> PROBE<1753> PROBE<1754> PROBE<1755> PROBE<1756> PROBE<1757>
+  PROBE<1758> PROBE<1759> PROBE<1760> PROBE<1761> PROBE<1762> PROBE<1763>
+  PROBE<1764> PROBE<1765> PROBE<1766> PROBE<1767> PROBE<1768> PROBE<1769>
+  PROBE<1770> PROBE<1771> PROBE<1772> PROBE<1773> PROBE<1774> PROBE<1775>
+  PROBE<1776> PROBE<1777> PROBE<1778> PROBE<1779> PROBE<1780> PROBE<1781>
+  PROBE<1782> PROBE<1783> PROBE<1784> PROBE<1785> PROBE<1786> PROBE<1787>
+  PROBE<1788> PROBE<1789> PROBE<1790> PROBE<1791> PROBE<1792> PROBE<1793>
+  PROBE<1794> PROBE<1795> PROBE<1796> PROBE<1797> PROBE<1798> PROBE<1799>
+  PROBE<1800> PROBE<1801> PROBE<1802> PROBE<1803> PROBE<1804> PROBE<1805>
+  PROBE<1806> PROBE<1807> PROBE<1808> PROBE<1809> PROBE<1810> PROBE<1811>
+  PROBE<1812> PROBE<1813> PROBE<1814> PROBE<1815> PROBE<1816> PROBE<1817>
+  PROBE<1818> PROBE<1819> PROBE<1820> PROBE<1821> PROBE<1822> PROBE<1823>
+  PROBE<1824> PROBE<1825> PROBE<1826> PROBE<1827> PROBE<1828> PROBE<1829>
+  PROBE<1830> PROBE<1831> PROBE<1832> PROBE<1833> PROBE<1834> PROBE<1835>
+  PROBE<1836> PROBE<1837> PROBE<1838> PROBE<1839> PROBE<1840> PROBE<1841>
+  PROBE<1842> PROBE<1843> PROBE<1844> PROBE<1845> PROBE<1846> PROBE<1847>
+  PROBE<1848> PROBE<1849> PROBE<1850> PROBE<1851> PROBE<1852> PROBE<1853>
+  PROBE<1854> PROBE<1855> PROBE<1856> PROBE<1857> PROBE<1858> PROBE<1859>
+  PROBE<1860> PROBE<1861> PROBE<1862> PROBE<1863> PROBE<1864> PROBE<1865>
+  PROBE<1866> PROBE<1867> PROBE<1868> PROBE<1869> PROBE<1870> PROBE<1871>
+  PROBE<1872> PROBE<1873> PROBE<1874> PROBE<1875> PROBE<1876> PROBE<1877>
+  PROBE<1878> PROBE<1879> PROBE<1880> PROBE<1881> PROBE<1882> PROBE<1883>
+  PROBE<1884> PROBE<1885> PROBE<1886> PROBE<1887> PROBE<1888> VDD VSS
* Connection: SBUS1, Terminal: CC_N_G_CC, Connection Key: ON
V479_to_CC_N_G_CC PROBE<479> VDD 0
V480_to_CC_N_G_CC PROBE<480> VDD 0
* Connection: SBUS1, Terminal: CC_P_G_CC, Connection Key: ON
V1427_to_CC_P_G_CC PROBE<1427> VDD 0
V1428_to_CC_P_G_CC PROBE<1428> VDD 0
* Connection: SBUS2, Terminal: CC_N_D_CC, Connection Key: ON
V531_to_CC_N_D_CC PROBE<531> VDD 0
V532_to_CC_N_D_CC PROBE<532> VDD 0
* Connection: SBUS2, Terminal: CC_P_D_CC, Connection Key: ON
V1479_to_CC_P_D_CC PROBE<1479> VDD 0
V1480_to_CC_P_D_CC PROBE<1480> VDD 0
* Connection: SBUS2, Terminal: DINV1_INP_L, Connection Key: ON
V55_to_DINV1_INP_L PROBE<55> VDD 0
V56_to_DINV1_INP_L PROBE<56> VDD 0
* Connection: SBUS2, Terminal: DINV1_INN_L, Connection Key: ON
V57_to_DINV1_INN_L PROBE<57> VDD 0
V58_to_DINV1_INN_L PROBE<58> VDD 0
* Connection: SBUS3, Terminal: DINV1_OUT_L, Connection Key: ON
V107_to_DINV1_OUT_L PROBE<107> VDD 0
V108_to_DINV1_OUT_L PROBE<108> VDD 0
* Connection: SBUS3, Terminal: DINV1_INP_R, Connection Key: ON
V109_to_DINV1_INP_R PROBE<109> VDD 0
V110_to_DINV1_INP_R PROBE<110> VDD 0
* Connection: SBUS3, Terminal: DINV1_INN_R, Connection Key: ON
V111_to_DINV1_INN_R PROBE<111> VDD 0
V112_to_DINV1_INN_R PROBE<112> VDD 0
* Connection: SBUS4, Terminal: DINV1_OUT_R, Connection Key: ON
V161_to_DINV1_OUT_R PROBE<161> VDD 0
V162_to_DINV1_OUT_R PROBE<162> VDD 0
* Connection: SBUS4, Terminal: DINV2_INP_L, Connection Key: ON
V163_to_DINV2_INP_L PROBE<163> VDD 0
V164_to_DINV2_INP_L PROBE<164> VDD 0
* Connection: SBUS4, Terminal: DINV2_INN_L, Connection Key: ON
V165_to_DINV2_INN_L PROBE<165> VDD 0
V166_to_DINV2_INN_L PROBE<166> VDD 0
* Connection: SBUS5, Terminal: DINV2_OUT_L, Connection Key: ON
V215_to_DINV2_OUT_L PROBE<215> VDD 0
V216_to_DINV2_OUT_L PROBE<216> VDD 0
* Connection: SBUS5, Terminal: DINV2_INP_R, Connection Key: ON
V217_to_DINV2_INP_R PROBE<217> VDD 0
V218_to_DINV2_INP_R PROBE<218> VDD 0
* Connection: SBUS5, Terminal: DINV2_INN_R, Connection Key: ON
V219_to_DINV2_INN_R PROBE<219> VDD 0
V220_to_DINV2_INN_R PROBE<220> VDD 0
* Connection: SBUS6, Terminal: DINV2_OUT_R, Connection Key: ON
V269_to_DINV2_OUT_R PROBE<269> VDD 0
V270_to_DINV2_OUT_R PROBE<270> VDD 0
* Connection: SBUS6, Terminal: DCC1_N_G_L_CC, Connection Key: ON
V1201_to_DCC1_N_G_L_CC PROBE<1201> VDD 0
V1202_to_DCC1_N_G_L_CC PROBE<1202> VDD 0
* Connection: SBUS6, Terminal: DCC1_P_G_L_CC, Connection Key: ON
V1691_to_DCC1_P_G_L_CC PROBE<1691> VDD 0
V1692_to_DCC1_P_G_L_CC PROBE<1692> VDD 0
* Connection: RBUS1, Pin: DCC1_N_D_L_CC, sw_matrix_pin: 59.0, Register: 1245
VDCC1_N_D_L_CC_to_RBUS1 PROBE<1245> VDD 0
* Connection: RBUS1, Pin: DCC1_P_D_L_CC, sw_matrix_pin: 1.0, Register: 289
VDCC1_P_D_L_CC_to_RBUS1 PROBE<289> VDD 0
* Connection: RBUS1, Pin: DCC1_N_G_R_CC, sw_matrix_pin: 57.0, Register: 1243
VDCC1_N_G_R_CC_to_RBUS1 PROBE<1243> VDD 0
* Connection: RBUS1, Pin: DCC1_P_G_R_CC, sw_matrix_pin: 89.0, Register: 1724
VDCC1_P_G_R_CC_to_RBUS1 PROBE<1724> VDD 0
* Connection: RBUS2, Pin: DCC1_N_D_R_CC, sw_matrix_pin: 61.0, Register: 1270
VDCC1_N_D_R_CC_to_RBUS2 PROBE<1270> VDD 0
* Connection: RBUS2, Pin: DCC1_P_D_R_CC, sw_matrix_pin: 3.0, Register: 314
VDCC1_P_D_R_CC_to_RBUS2 PROBE<314> VDD 0
* Connection: RBUS2, Pin: DCC2_N_G_L_CC, sw_matrix_pin: 31.0, Register: 791
VDCC2_N_G_L_CC_to_RBUS2 PROBE<791> VDD 0
* Connection: RBUS2, Pin: DCC2_P_G_L_CC, sw_matrix_pin: 64.0, Register: 1273
VDCC2_P_G_L_CC_to_RBUS2 PROBE<1273> VDD 0
* Connection: RBUS3, Pin: DCC2_N_D_L_CC, sw_matrix_pin: 35.0, Register: 818
VDCC2_N_D_L_CC_to_RBUS3 PROBE<818> VDD 0
* Connection: RBUS3, Pin: DCC2_P_D_L_CC, sw_matrix_pin: 68.0, Register: 1300
VDCC2_P_D_L_CC_to_RBUS3 PROBE<1300> VDD 0
* Connection: RBUS3, Pin: DCC2_N_G_R_CC, sw_matrix_pin: 33.0, Register: 816
VDCC2_N_G_R_CC_to_RBUS3 PROBE<816> VDD 0
* Connection: RBUS3, Pin: DCC2_P_G_R_CC, sw_matrix_pin: 66.0, Register: 1298
VDCC2_P_G_R_CC_to_RBUS3 PROBE<1298> VDD 0
* Connection: RBUS4, Pin: DCC2_N_D_R_CC, sw_matrix_pin: 37.0, Register: 843
VDCC2_N_D_R_CC_to_RBUS4 PROBE<843> VDD 0
* Connection: RBUS4, Pin: DCC2_P_D_R_CC, sw_matrix_pin: 70.0, Register: 1774
VDCC2_P_D_R_CC_to_RBUS4 PROBE<1774> VDD 0
* Connection: RBUS4, Pin: DCC3_N_G_L_CC, sw_matrix_pin: 39.0, Register: 845
VDCC3_N_G_L_CC_to_RBUS4 PROBE<845> VDD 0
* Connection: RBUS4, Pin: DCC3_P_G_L_CC, sw_matrix_pin: 48.0, Register: 1303
VDCC3_P_G_L_CC_to_RBUS4 PROBE<1303> VDD 0
* Connection: RBUS5, Pin: DCC3_N_D_L_CC, sw_matrix_pin: 43.0, Register: 872
VDCC3_N_D_L_CC_to_RBUS5 PROBE<872> VDD 0
* Connection: RBUS5, Pin: DCC3_P_D_L_CC, sw_matrix_pin: 52.0, Register: 1330
VDCC3_P_D_L_CC_to_RBUS5 PROBE<1330> VDD 0
* Connection: RBUS5, Pin: DCC3_N_G_R_CC, sw_matrix_pin: 41.0, Register: 870
VDCC3_N_G_R_CC_to_RBUS5 PROBE<870> VDD 0
* Connection: RBUS5, Pin: DCC3_P_G_R_CC, sw_matrix_pin: 50.0, Register: 1328
VDCC3_P_G_R_CC_to_RBUS5 PROBE<1328> VDD 0
* Connection: RBUS8, Pin: VDD, sw_matrix_pin: 91.0, Register: 1887
VVDD_to_RBUS8 PROBE<1887> VDD 0
* Connection: RBUS8, Pin: CC_N_G_CS, sw_matrix_pin: 28.0, Register: 926
VCC_N_G_CS_to_RBUS8 PROBE<926> VDD 0
* Connection: RBUS8, Pin: DCC1_N_G_L_CS, sw_matrix_pin: 56.0, Register: 1403
VDCC1_N_G_L_CS_to_RBUS8 PROBE<1403> VDD 0
* Connection: RBUS8, Pin: DCC1_N_G_R_CS, sw_matrix_pin: 58.0, Register: 1405
VDCC1_N_G_R_CS_to_RBUS8 PROBE<1405> VDD 0
* Connection: RBUS8, Pin: DCC2_N_G_L_CS, sw_matrix_pin: 32.0, Register: 930
VDCC2_N_G_L_CS_to_RBUS8 PROBE<930> VDD 0
* Connection: RBUS8, Pin: DCC2_N_G_R_CS, sw_matrix_pin: 34.0, Register: 932
VDCC2_N_G_R_CS_to_RBUS8 PROBE<932> VDD 0
* Connection: RBUS8, Pin: DCC3_N_G_L_CS, sw_matrix_pin: 40.0, Register: 938
VDCC3_N_G_L_CS_to_RBUS8 PROBE<938> VDD 0
* Connection: RBUS8, Pin: DCC3_N_G_R_CS, sw_matrix_pin: 42.0, Register: 940
VDCC3_N_G_R_CS_to_RBUS8 PROBE<940> VDD 0
* Connection: RBUS8, Pin: DCC4_P_G_L_CS, sw_matrix_pin: 17.0, Register: 466
VDCC4_P_G_L_CS_to_RBUS8 PROBE<466> VDD 0
* Connection: RBUS8, Pin: DCC4_P_G_R_CS, sw_matrix_pin: 19.0, Register: 468
VDCC4_P_G_R_CS_to_RBUS8 PROBE<468> VDD 0
* Connection: RBUS7, Pin: VSS, sw_matrix_pin: 92.0, Register: 1865
VVSS_to_RBUS7 PROBE<1865> VDD 0
* Connection: RBUS7, Pin: CC_P_G_CS, sw_matrix_pin: 74.0, Register: 1847
VCC_P_G_CS_to_RBUS7 PROBE<1847> VDD 0
* Connection: RBUS7, Pin: DCC1_P_G_L_CS, sw_matrix_pin: 86.0, Register: 1859
VDCC1_P_G_L_CS_to_RBUS7 PROBE<1859> VDD 0
* Connection: RBUS7, Pin: DCC1_P_G_R_CS, sw_matrix_pin: 88.0, Register: 1861
VDCC1_P_G_R_CS_to_RBUS7 PROBE<1861> VDD 0
* Connection: RBUS7, Pin: DCC2_P_G_L_CS, sw_matrix_pin: 63.0, Register: 1387
VDCC2_P_G_L_CS_to_RBUS7 PROBE<1387> VDD 0
* Connection: RBUS7, Pin: DCC2_P_G_R_CS, sw_matrix_pin: 65.0, Register: 1389
VDCC2_P_G_R_CS_to_RBUS7 PROBE<1389> VDD 0
* Connection: RBUS7, Pin: DCC3_P_G_L_CS, sw_matrix_pin: 47.0, Register: 1371
VDCC3_P_G_L_CS_to_RBUS7 PROBE<1371> VDD 0
* Connection: RBUS7, Pin: DCC3_P_G_R_CS, sw_matrix_pin: 49.0, Register: 1373
VDCC3_P_G_R_CS_to_RBUS7 PROBE<1373> VDD 0
* Connection: RBUS7, Pin: DCC4_N_G_L_CS, sw_matrix_pin: 79.0, Register: 1852
VDCC4_N_G_L_CS_to_RBUS7 PROBE<1852> VDD 0
* Connection: RBUS7, Pin: DCC4_N_G_R_CS, sw_matrix_pin: 81.0, Register: 1854
VDCC4_N_G_R_CS_to_RBUS7 PROBE<1854> VDD 0
Vprobe_1_to_VSS PROBE<1> VSS 0
Vprobe_2_to_VSS PROBE<2> VSS 0
Vprobe_3_to_VSS PROBE<3> VSS 0
Vprobe_4_to_VSS PROBE<4> VSS 0
Vprobe_5_to_VSS PROBE<5> VSS 0
Vprobe_6_to_VSS PROBE<6> VSS 0
Vprobe_7_to_VSS PROBE<7> VSS 0
Vprobe_8_to_VSS PROBE<8> VSS 0
Vprobe_9_to_VSS PROBE<9> VSS 0
Vprobe_10_to_VSS PROBE<10> VSS 0
Vprobe_11_to_VSS PROBE<11> VSS 0
Vprobe_12_to_VSS PROBE<12> VSS 0
Vprobe_13_to_VSS PROBE<13> VSS 0
Vprobe_14_to_VSS PROBE<14> VSS 0
Vprobe_15_to_VSS PROBE<15> VSS 0
Vprobe_16_to_VSS PROBE<16> VSS 0
Vprobe_17_to_VSS PROBE<17> VSS 0
Vprobe_18_to_VSS PROBE<18> VSS 0
Vprobe_19_to_VSS PROBE<19> VSS 0
Vprobe_20_to_VSS PROBE<20> VSS 0
Vprobe_21_to_VSS PROBE<21> VSS 0
Vprobe_22_to_VSS PROBE<22> VSS 0
Vprobe_23_to_VSS PROBE<23> VSS 0
Vprobe_24_to_VSS PROBE<24> VSS 0
Vprobe_25_to_VSS PROBE<25> VSS 0
Vprobe_26_to_VSS PROBE<26> VSS 0
Vprobe_27_to_VSS PROBE<27> VSS 0
Vprobe_28_to_VSS PROBE<28> VSS 0
Vprobe_29_to_VSS PROBE<29> VSS 0
Vprobe_30_to_VSS PROBE<30> VSS 0
Vprobe_31_to_VSS PROBE<31> VSS 0
Vprobe_32_to_VSS PROBE<32> VSS 0
Vprobe_33_to_VSS PROBE<33> VSS 0
Vprobe_34_to_VSS PROBE<34> VSS 0
Vprobe_35_to_VSS PROBE<35> VSS 0
Vprobe_36_to_VSS PROBE<36> VSS 0
Vprobe_37_to_VSS PROBE<37> VSS 0
Vprobe_38_to_VSS PROBE<38> VSS 0
Vprobe_39_to_VSS PROBE<39> VSS 0
Vprobe_40_to_VSS PROBE<40> VSS 0
Vprobe_41_to_VSS PROBE<41> VSS 0
Vprobe_42_to_VSS PROBE<42> VSS 0
Vprobe_43_to_VSS PROBE<43> VSS 0
Vprobe_44_to_VSS PROBE<44> VSS 0
Vprobe_45_to_VSS PROBE<45> VSS 0
Vprobe_46_to_VSS PROBE<46> VSS 0
Vprobe_47_to_VSS PROBE<47> VSS 0
Vprobe_48_to_VSS PROBE<48> VSS 0
Vprobe_49_to_VSS PROBE<49> VSS 0
Vprobe_50_to_VSS PROBE<50> VSS 0
Vprobe_51_to_VSS PROBE<51> VSS 0
Vprobe_52_to_VSS PROBE<52> VSS 0
Vprobe_53_to_VSS PROBE<53> VSS 0
Vprobe_54_to_VSS PROBE<54> VSS 0
Vprobe_59_to_VSS PROBE<59> VSS 0
Vprobe_60_to_VSS PROBE<60> VSS 0
Vprobe_61_to_VSS PROBE<61> VSS 0
Vprobe_62_to_VSS PROBE<62> VSS 0
Vprobe_63_to_VSS PROBE<63> VSS 0
Vprobe_64_to_VSS PROBE<64> VSS 0
Vprobe_65_to_VSS PROBE<65> VSS 0
Vprobe_66_to_VSS PROBE<66> VSS 0
Vprobe_67_to_VSS PROBE<67> VSS 0
Vprobe_68_to_VSS PROBE<68> VSS 0
Vprobe_69_to_VSS PROBE<69> VSS 0
Vprobe_70_to_VSS PROBE<70> VSS 0
Vprobe_71_to_VSS PROBE<71> VSS 0
Vprobe_72_to_VSS PROBE<72> VSS 0
Vprobe_73_to_VSS PROBE<73> VSS 0
Vprobe_74_to_VSS PROBE<74> VSS 0
Vprobe_75_to_VSS PROBE<75> VSS 0
Vprobe_76_to_VSS PROBE<76> VSS 0
Vprobe_77_to_VSS PROBE<77> VSS 0
Vprobe_78_to_VSS PROBE<78> VSS 0
Vprobe_79_to_VSS PROBE<79> VSS 0
Vprobe_80_to_VSS PROBE<80> VSS 0
Vprobe_81_to_VSS PROBE<81> VSS 0
Vprobe_82_to_VSS PROBE<82> VSS 0
Vprobe_83_to_VSS PROBE<83> VSS 0
Vprobe_84_to_VSS PROBE<84> VSS 0
Vprobe_85_to_VSS PROBE<85> VSS 0
Vprobe_86_to_VSS PROBE<86> VSS 0
Vprobe_87_to_VSS PROBE<87> VSS 0
Vprobe_88_to_VSS PROBE<88> VSS 0
Vprobe_89_to_VSS PROBE<89> VSS 0
Vprobe_90_to_VSS PROBE<90> VSS 0
Vprobe_91_to_VSS PROBE<91> VSS 0
Vprobe_92_to_VSS PROBE<92> VSS 0
Vprobe_93_to_VSS PROBE<93> VSS 0
Vprobe_94_to_VSS PROBE<94> VSS 0
Vprobe_95_to_VSS PROBE<95> VSS 0
Vprobe_96_to_VSS PROBE<96> VSS 0
Vprobe_97_to_VSS PROBE<97> VSS 0
Vprobe_98_to_VSS PROBE<98> VSS 0
Vprobe_99_to_VSS PROBE<99> VSS 0
Vprobe_100_to_VSS PROBE<100> VSS 0
Vprobe_101_to_VSS PROBE<101> VSS 0
Vprobe_102_to_VSS PROBE<102> VSS 0
Vprobe_103_to_VSS PROBE<103> VSS 0
Vprobe_104_to_VSS PROBE<104> VSS 0
Vprobe_105_to_VSS PROBE<105> VSS 0
Vprobe_106_to_VSS PROBE<106> VSS 0
Vprobe_113_to_VSS PROBE<113> VSS 0
Vprobe_114_to_VSS PROBE<114> VSS 0
Vprobe_115_to_VSS PROBE<115> VSS 0
Vprobe_116_to_VSS PROBE<116> VSS 0
Vprobe_117_to_VSS PROBE<117> VSS 0
Vprobe_118_to_VSS PROBE<118> VSS 0
Vprobe_119_to_VSS PROBE<119> VSS 0
Vprobe_120_to_VSS PROBE<120> VSS 0
Vprobe_121_to_VSS PROBE<121> VSS 0
Vprobe_122_to_VSS PROBE<122> VSS 0
Vprobe_123_to_VSS PROBE<123> VSS 0
Vprobe_124_to_VSS PROBE<124> VSS 0
Vprobe_125_to_VSS PROBE<125> VSS 0
Vprobe_126_to_VSS PROBE<126> VSS 0
Vprobe_127_to_VSS PROBE<127> VSS 0
Vprobe_128_to_VSS PROBE<128> VSS 0
Vprobe_129_to_VSS PROBE<129> VSS 0
Vprobe_130_to_VSS PROBE<130> VSS 0
Vprobe_131_to_VSS PROBE<131> VSS 0
Vprobe_132_to_VSS PROBE<132> VSS 0
Vprobe_133_to_VSS PROBE<133> VSS 0
Vprobe_134_to_VSS PROBE<134> VSS 0
Vprobe_135_to_VSS PROBE<135> VSS 0
Vprobe_136_to_VSS PROBE<136> VSS 0
Vprobe_137_to_VSS PROBE<137> VSS 0
Vprobe_138_to_VSS PROBE<138> VSS 0
Vprobe_139_to_VSS PROBE<139> VSS 0
Vprobe_140_to_VSS PROBE<140> VSS 0
Vprobe_141_to_VSS PROBE<141> VSS 0
Vprobe_142_to_VSS PROBE<142> VSS 0
Vprobe_143_to_VSS PROBE<143> VSS 0
Vprobe_144_to_VSS PROBE<144> VSS 0
Vprobe_145_to_VSS PROBE<145> VSS 0
Vprobe_146_to_VSS PROBE<146> VSS 0
Vprobe_147_to_VSS PROBE<147> VSS 0
Vprobe_148_to_VSS PROBE<148> VSS 0
Vprobe_149_to_VSS PROBE<149> VSS 0
Vprobe_150_to_VSS PROBE<150> VSS 0
Vprobe_151_to_VSS PROBE<151> VSS 0
Vprobe_152_to_VSS PROBE<152> VSS 0
Vprobe_153_to_VSS PROBE<153> VSS 0
Vprobe_154_to_VSS PROBE<154> VSS 0
Vprobe_155_to_VSS PROBE<155> VSS 0
Vprobe_156_to_VSS PROBE<156> VSS 0
Vprobe_157_to_VSS PROBE<157> VSS 0
Vprobe_158_to_VSS PROBE<158> VSS 0
Vprobe_159_to_VSS PROBE<159> VSS 0
Vprobe_160_to_VSS PROBE<160> VSS 0
Vprobe_167_to_VSS PROBE<167> VSS 0
Vprobe_168_to_VSS PROBE<168> VSS 0
Vprobe_169_to_VSS PROBE<169> VSS 0
Vprobe_170_to_VSS PROBE<170> VSS 0
Vprobe_171_to_VSS PROBE<171> VSS 0
Vprobe_172_to_VSS PROBE<172> VSS 0
Vprobe_173_to_VSS PROBE<173> VSS 0
Vprobe_174_to_VSS PROBE<174> VSS 0
Vprobe_175_to_VSS PROBE<175> VSS 0
Vprobe_176_to_VSS PROBE<176> VSS 0
Vprobe_177_to_VSS PROBE<177> VSS 0
Vprobe_178_to_VSS PROBE<178> VSS 0
Vprobe_179_to_VSS PROBE<179> VSS 0
Vprobe_180_to_VSS PROBE<180> VSS 0
Vprobe_181_to_VSS PROBE<181> VSS 0
Vprobe_182_to_VSS PROBE<182> VSS 0
Vprobe_183_to_VSS PROBE<183> VSS 0
Vprobe_184_to_VSS PROBE<184> VSS 0
Vprobe_185_to_VSS PROBE<185> VSS 0
Vprobe_186_to_VSS PROBE<186> VSS 0
Vprobe_187_to_VSS PROBE<187> VSS 0
Vprobe_188_to_VSS PROBE<188> VSS 0
Vprobe_189_to_VSS PROBE<189> VSS 0
Vprobe_190_to_VSS PROBE<190> VSS 0
Vprobe_191_to_VSS PROBE<191> VSS 0
Vprobe_192_to_VSS PROBE<192> VSS 0
Vprobe_193_to_VSS PROBE<193> VSS 0
Vprobe_194_to_VSS PROBE<194> VSS 0
Vprobe_195_to_VSS PROBE<195> VSS 0
Vprobe_196_to_VSS PROBE<196> VSS 0
Vprobe_197_to_VSS PROBE<197> VSS 0
Vprobe_198_to_VSS PROBE<198> VSS 0
Vprobe_199_to_VSS PROBE<199> VSS 0
Vprobe_200_to_VSS PROBE<200> VSS 0
Vprobe_201_to_VSS PROBE<201> VSS 0
Vprobe_202_to_VSS PROBE<202> VSS 0
Vprobe_203_to_VSS PROBE<203> VSS 0
Vprobe_204_to_VSS PROBE<204> VSS 0
Vprobe_205_to_VSS PROBE<205> VSS 0
Vprobe_206_to_VSS PROBE<206> VSS 0
Vprobe_207_to_VSS PROBE<207> VSS 0
Vprobe_208_to_VSS PROBE<208> VSS 0
Vprobe_209_to_VSS PROBE<209> VSS 0
Vprobe_210_to_VSS PROBE<210> VSS 0
Vprobe_211_to_VSS PROBE<211> VSS 0
Vprobe_212_to_VSS PROBE<212> VSS 0
Vprobe_213_to_VSS PROBE<213> VSS 0
Vprobe_214_to_VSS PROBE<214> VSS 0
Vprobe_221_to_VSS PROBE<221> VSS 0
Vprobe_222_to_VSS PROBE<222> VSS 0
Vprobe_223_to_VSS PROBE<223> VSS 0
Vprobe_224_to_VSS PROBE<224> VSS 0
Vprobe_225_to_VSS PROBE<225> VSS 0
Vprobe_226_to_VSS PROBE<226> VSS 0
Vprobe_227_to_VSS PROBE<227> VSS 0
Vprobe_228_to_VSS PROBE<228> VSS 0
Vprobe_229_to_VSS PROBE<229> VSS 0
Vprobe_230_to_VSS PROBE<230> VSS 0
Vprobe_231_to_VSS PROBE<231> VSS 0
Vprobe_232_to_VSS PROBE<232> VSS 0
Vprobe_233_to_VSS PROBE<233> VSS 0
Vprobe_234_to_VSS PROBE<234> VSS 0
Vprobe_235_to_VSS PROBE<235> VSS 0
Vprobe_236_to_VSS PROBE<236> VSS 0
Vprobe_237_to_VSS PROBE<237> VSS 0
Vprobe_238_to_VSS PROBE<238> VSS 0
Vprobe_239_to_VSS PROBE<239> VSS 0
Vprobe_240_to_VSS PROBE<240> VSS 0
Vprobe_241_to_VSS PROBE<241> VSS 0
Vprobe_242_to_VSS PROBE<242> VSS 0
Vprobe_243_to_VSS PROBE<243> VSS 0
Vprobe_244_to_VSS PROBE<244> VSS 0
Vprobe_245_to_VSS PROBE<245> VSS 0
Vprobe_246_to_VSS PROBE<246> VSS 0
Vprobe_247_to_VSS PROBE<247> VSS 0
Vprobe_248_to_VSS PROBE<248> VSS 0
Vprobe_249_to_VSS PROBE<249> VSS 0
Vprobe_250_to_VSS PROBE<250> VSS 0
Vprobe_251_to_VSS PROBE<251> VSS 0
Vprobe_252_to_VSS PROBE<252> VSS 0
Vprobe_253_to_VSS PROBE<253> VSS 0
Vprobe_254_to_VSS PROBE<254> VSS 0
Vprobe_255_to_VSS PROBE<255> VSS 0
Vprobe_256_to_VSS PROBE<256> VSS 0
Vprobe_257_to_VSS PROBE<257> VSS 0
Vprobe_258_to_VSS PROBE<258> VSS 0
Vprobe_259_to_VSS PROBE<259> VSS 0
Vprobe_260_to_VSS PROBE<260> VSS 0
Vprobe_261_to_VSS PROBE<261> VSS 0
Vprobe_262_to_VSS PROBE<262> VSS 0
Vprobe_263_to_VSS PROBE<263> VSS 0
Vprobe_264_to_VSS PROBE<264> VSS 0
Vprobe_265_to_VSS PROBE<265> VSS 0
Vprobe_266_to_VSS PROBE<266> VSS 0
Vprobe_267_to_VSS PROBE<267> VSS 0
Vprobe_268_to_VSS PROBE<268> VSS 0
Vprobe_271_to_VSS PROBE<271> VSS 0
Vprobe_272_to_VSS PROBE<272> VSS 0
Vprobe_273_to_VSS PROBE<273> VSS 0
Vprobe_274_to_VSS PROBE<274> VSS 0
Vprobe_275_to_VSS PROBE<275> VSS 0
Vprobe_276_to_VSS PROBE<276> VSS 0
Vprobe_277_to_VSS PROBE<277> VSS 0
Vprobe_278_to_VSS PROBE<278> VSS 0
Vprobe_279_to_VSS PROBE<279> VSS 0
Vprobe_280_to_VSS PROBE<280> VSS 0
Vprobe_281_to_VSS PROBE<281> VSS 0
Vprobe_282_to_VSS PROBE<282> VSS 0
Vprobe_283_to_VSS PROBE<283> VSS 0
Vprobe_284_to_VSS PROBE<284> VSS 0
Vprobe_285_to_VSS PROBE<285> VSS 0
Vprobe_286_to_VSS PROBE<286> VSS 0
Vprobe_287_to_VSS PROBE<287> VSS 0
Vprobe_288_to_VSS PROBE<288> VSS 0
Vprobe_290_to_VSS PROBE<290> VSS 0
Vprobe_291_to_VSS PROBE<291> VSS 0
Vprobe_292_to_VSS PROBE<292> VSS 0
Vprobe_293_to_VSS PROBE<293> VSS 0
Vprobe_294_to_VSS PROBE<294> VSS 0
Vprobe_295_to_VSS PROBE<295> VSS 0
Vprobe_296_to_VSS PROBE<296> VSS 0
Vprobe_297_to_VSS PROBE<297> VSS 0
Vprobe_298_to_VSS PROBE<298> VSS 0
Vprobe_299_to_VSS PROBE<299> VSS 0
Vprobe_300_to_VSS PROBE<300> VSS 0
Vprobe_301_to_VSS PROBE<301> VSS 0
Vprobe_302_to_VSS PROBE<302> VSS 0
Vprobe_303_to_VSS PROBE<303> VSS 0
Vprobe_304_to_VSS PROBE<304> VSS 0
Vprobe_305_to_VSS PROBE<305> VSS 0
Vprobe_306_to_VSS PROBE<306> VSS 0
Vprobe_307_to_VSS PROBE<307> VSS 0
Vprobe_308_to_VSS PROBE<308> VSS 0
Vprobe_309_to_VSS PROBE<309> VSS 0
Vprobe_310_to_VSS PROBE<310> VSS 0
Vprobe_311_to_VSS PROBE<311> VSS 0
Vprobe_312_to_VSS PROBE<312> VSS 0
Vprobe_313_to_VSS PROBE<313> VSS 0
Vprobe_315_to_VSS PROBE<315> VSS 0
Vprobe_316_to_VSS PROBE<316> VSS 0
Vprobe_317_to_VSS PROBE<317> VSS 0
Vprobe_318_to_VSS PROBE<318> VSS 0
Vprobe_319_to_VSS PROBE<319> VSS 0
Vprobe_320_to_VSS PROBE<320> VSS 0
Vprobe_321_to_VSS PROBE<321> VSS 0
Vprobe_322_to_VSS PROBE<322> VSS 0
Vprobe_323_to_VSS PROBE<323> VSS 0
Vprobe_324_to_VSS PROBE<324> VSS 0
Vprobe_325_to_VSS PROBE<325> VSS 0
Vprobe_326_to_VSS PROBE<326> VSS 0
Vprobe_327_to_VSS PROBE<327> VSS 0
Vprobe_328_to_VSS PROBE<328> VSS 0
Vprobe_329_to_VSS PROBE<329> VSS 0
Vprobe_330_to_VSS PROBE<330> VSS 0
Vprobe_331_to_VSS PROBE<331> VSS 0
Vprobe_332_to_VSS PROBE<332> VSS 0
Vprobe_333_to_VSS PROBE<333> VSS 0
Vprobe_334_to_VSS PROBE<334> VSS 0
Vprobe_335_to_VSS PROBE<335> VSS 0
Vprobe_336_to_VSS PROBE<336> VSS 0
Vprobe_337_to_VSS PROBE<337> VSS 0
Vprobe_338_to_VSS PROBE<338> VSS 0
Vprobe_339_to_VSS PROBE<339> VSS 0
Vprobe_340_to_VSS PROBE<340> VSS 0
Vprobe_341_to_VSS PROBE<341> VSS 0
Vprobe_342_to_VSS PROBE<342> VSS 0
Vprobe_343_to_VSS PROBE<343> VSS 0
Vprobe_344_to_VSS PROBE<344> VSS 0
Vprobe_345_to_VSS PROBE<345> VSS 0
Vprobe_346_to_VSS PROBE<346> VSS 0
Vprobe_347_to_VSS PROBE<347> VSS 0
Vprobe_348_to_VSS PROBE<348> VSS 0
Vprobe_349_to_VSS PROBE<349> VSS 0
Vprobe_350_to_VSS PROBE<350> VSS 0
Vprobe_351_to_VSS PROBE<351> VSS 0
Vprobe_352_to_VSS PROBE<352> VSS 0
Vprobe_353_to_VSS PROBE<353> VSS 0
Vprobe_354_to_VSS PROBE<354> VSS 0
Vprobe_355_to_VSS PROBE<355> VSS 0
Vprobe_356_to_VSS PROBE<356> VSS 0
Vprobe_357_to_VSS PROBE<357> VSS 0
Vprobe_358_to_VSS PROBE<358> VSS 0
Vprobe_359_to_VSS PROBE<359> VSS 0
Vprobe_360_to_VSS PROBE<360> VSS 0
Vprobe_361_to_VSS PROBE<361> VSS 0
Vprobe_362_to_VSS PROBE<362> VSS 0
Vprobe_363_to_VSS PROBE<363> VSS 0
Vprobe_364_to_VSS PROBE<364> VSS 0
Vprobe_365_to_VSS PROBE<365> VSS 0
Vprobe_366_to_VSS PROBE<366> VSS 0
Vprobe_367_to_VSS PROBE<367> VSS 0
Vprobe_368_to_VSS PROBE<368> VSS 0
Vprobe_369_to_VSS PROBE<369> VSS 0
Vprobe_370_to_VSS PROBE<370> VSS 0
Vprobe_371_to_VSS PROBE<371> VSS 0
Vprobe_372_to_VSS PROBE<372> VSS 0
Vprobe_373_to_VSS PROBE<373> VSS 0
Vprobe_374_to_VSS PROBE<374> VSS 0
Vprobe_375_to_VSS PROBE<375> VSS 0
Vprobe_376_to_VSS PROBE<376> VSS 0
Vprobe_377_to_VSS PROBE<377> VSS 0
Vprobe_378_to_VSS PROBE<378> VSS 0
Vprobe_379_to_VSS PROBE<379> VSS 0
Vprobe_380_to_VSS PROBE<380> VSS 0
Vprobe_381_to_VSS PROBE<381> VSS 0
Vprobe_382_to_VSS PROBE<382> VSS 0
Vprobe_383_to_VSS PROBE<383> VSS 0
Vprobe_384_to_VSS PROBE<384> VSS 0
Vprobe_385_to_VSS PROBE<385> VSS 0
Vprobe_386_to_VSS PROBE<386> VSS 0
Vprobe_387_to_VSS PROBE<387> VSS 0
Vprobe_388_to_VSS PROBE<388> VSS 0
Vprobe_389_to_VSS PROBE<389> VSS 0
Vprobe_390_to_VSS PROBE<390> VSS 0
Vprobe_391_to_VSS PROBE<391> VSS 0
Vprobe_392_to_VSS PROBE<392> VSS 0
Vprobe_393_to_VSS PROBE<393> VSS 0
Vprobe_394_to_VSS PROBE<394> VSS 0
Vprobe_395_to_VSS PROBE<395> VSS 0
Vprobe_396_to_VSS PROBE<396> VSS 0
Vprobe_397_to_VSS PROBE<397> VSS 0
Vprobe_398_to_VSS PROBE<398> VSS 0
Vprobe_399_to_VSS PROBE<399> VSS 0
Vprobe_400_to_VSS PROBE<400> VSS 0
Vprobe_401_to_VSS PROBE<401> VSS 0
Vprobe_402_to_VSS PROBE<402> VSS 0
Vprobe_403_to_VSS PROBE<403> VSS 0
Vprobe_404_to_VSS PROBE<404> VSS 0
Vprobe_405_to_VSS PROBE<405> VSS 0
Vprobe_406_to_VSS PROBE<406> VSS 0
Vprobe_407_to_VSS PROBE<407> VSS 0
Vprobe_408_to_VSS PROBE<408> VSS 0
Vprobe_409_to_VSS PROBE<409> VSS 0
Vprobe_410_to_VSS PROBE<410> VSS 0
Vprobe_411_to_VSS PROBE<411> VSS 0
Vprobe_412_to_VSS PROBE<412> VSS 0
Vprobe_413_to_VSS PROBE<413> VSS 0
Vprobe_414_to_VSS PROBE<414> VSS 0
Vprobe_415_to_VSS PROBE<415> VSS 0
Vprobe_416_to_VSS PROBE<416> VSS 0
Vprobe_417_to_VSS PROBE<417> VSS 0
Vprobe_418_to_VSS PROBE<418> VSS 0
Vprobe_419_to_VSS PROBE<419> VSS 0
Vprobe_420_to_VSS PROBE<420> VSS 0
Vprobe_421_to_VSS PROBE<421> VSS 0
Vprobe_422_to_VSS PROBE<422> VSS 0
Vprobe_423_to_VSS PROBE<423> VSS 0
Vprobe_424_to_VSS PROBE<424> VSS 0
Vprobe_425_to_VSS PROBE<425> VSS 0
Vprobe_426_to_VSS PROBE<426> VSS 0
Vprobe_427_to_VSS PROBE<427> VSS 0
Vprobe_428_to_VSS PROBE<428> VSS 0
Vprobe_429_to_VSS PROBE<429> VSS 0
Vprobe_430_to_VSS PROBE<430> VSS 0
Vprobe_431_to_VSS PROBE<431> VSS 0
Vprobe_432_to_VSS PROBE<432> VSS 0
Vprobe_433_to_VSS PROBE<433> VSS 0
Vprobe_434_to_VSS PROBE<434> VSS 0
Vprobe_435_to_VSS PROBE<435> VSS 0
Vprobe_436_to_VSS PROBE<436> VSS 0
Vprobe_437_to_VSS PROBE<437> VSS 0
Vprobe_438_to_VSS PROBE<438> VSS 0
Vprobe_439_to_VSS PROBE<439> VSS 0
Vprobe_440_to_VSS PROBE<440> VSS 0
Vprobe_441_to_VSS PROBE<441> VSS 0
Vprobe_442_to_VSS PROBE<442> VSS 0
Vprobe_443_to_VSS PROBE<443> VSS 0
Vprobe_444_to_VSS PROBE<444> VSS 0
Vprobe_445_to_VSS PROBE<445> VSS 0
Vprobe_446_to_VSS PROBE<446> VSS 0
Vprobe_447_to_VSS PROBE<447> VSS 0
Vprobe_448_to_VSS PROBE<448> VSS 0
Vprobe_449_to_VSS PROBE<449> VSS 0
Vprobe_450_to_VSS PROBE<450> VSS 0
Vprobe_451_to_VSS PROBE<451> VSS 0
Vprobe_452_to_VSS PROBE<452> VSS 0
Vprobe_453_to_VSS PROBE<453> VSS 0
Vprobe_454_to_VSS PROBE<454> VSS 0
Vprobe_455_to_VSS PROBE<455> VSS 0
Vprobe_456_to_VSS PROBE<456> VSS 0
Vprobe_457_to_VSS PROBE<457> VSS 0
Vprobe_458_to_VSS PROBE<458> VSS 0
Vprobe_459_to_VSS PROBE<459> VSS 0
Vprobe_460_to_VSS PROBE<460> VSS 0
Vprobe_461_to_VSS PROBE<461> VSS 0
Vprobe_462_to_VSS PROBE<462> VSS 0
Vprobe_463_to_VSS PROBE<463> VSS 0
Vprobe_464_to_VSS PROBE<464> VSS 0
Vprobe_465_to_VSS PROBE<465> VSS 0
Vprobe_467_to_VSS PROBE<467> VSS 0
Vprobe_469_to_VSS PROBE<469> VSS 0
Vprobe_470_to_VSS PROBE<470> VSS 0
Vprobe_471_to_VSS PROBE<471> VSS 0
Vprobe_472_to_VSS PROBE<472> VSS 0
Vprobe_473_to_VSS PROBE<473> VSS 0
Vprobe_474_to_VSS PROBE<474> VSS 0
Vprobe_475_to_VSS PROBE<475> VSS 0
Vprobe_476_to_VSS PROBE<476> VSS 0
Vprobe_477_to_VSS PROBE<477> VSS 0
Vprobe_478_to_VSS PROBE<478> VSS 0
Vprobe_481_to_VSS PROBE<481> VSS 0
Vprobe_482_to_VSS PROBE<482> VSS 0
Vprobe_483_to_VSS PROBE<483> VSS 0
Vprobe_484_to_VSS PROBE<484> VSS 0
Vprobe_485_to_VSS PROBE<485> VSS 0
Vprobe_486_to_VSS PROBE<486> VSS 0
Vprobe_487_to_VSS PROBE<487> VSS 0
Vprobe_488_to_VSS PROBE<488> VSS 0
Vprobe_489_to_VSS PROBE<489> VSS 0
Vprobe_490_to_VSS PROBE<490> VSS 0
Vprobe_491_to_VSS PROBE<491> VSS 0
Vprobe_492_to_VSS PROBE<492> VSS 0
Vprobe_493_to_VSS PROBE<493> VSS 0
Vprobe_494_to_VSS PROBE<494> VSS 0
Vprobe_495_to_VSS PROBE<495> VSS 0
Vprobe_496_to_VSS PROBE<496> VSS 0
Vprobe_497_to_VSS PROBE<497> VSS 0
Vprobe_498_to_VSS PROBE<498> VSS 0
Vprobe_499_to_VSS PROBE<499> VSS 0
Vprobe_500_to_VSS PROBE<500> VSS 0
Vprobe_501_to_VSS PROBE<501> VSS 0
Vprobe_502_to_VSS PROBE<502> VSS 0
Vprobe_503_to_VSS PROBE<503> VSS 0
Vprobe_504_to_VSS PROBE<504> VSS 0
Vprobe_505_to_VSS PROBE<505> VSS 0
Vprobe_506_to_VSS PROBE<506> VSS 0
Vprobe_507_to_VSS PROBE<507> VSS 0
Vprobe_508_to_VSS PROBE<508> VSS 0
Vprobe_509_to_VSS PROBE<509> VSS 0
Vprobe_510_to_VSS PROBE<510> VSS 0
Vprobe_511_to_VSS PROBE<511> VSS 0
Vprobe_512_to_VSS PROBE<512> VSS 0
Vprobe_513_to_VSS PROBE<513> VSS 0
Vprobe_514_to_VSS PROBE<514> VSS 0
Vprobe_515_to_VSS PROBE<515> VSS 0
Vprobe_516_to_VSS PROBE<516> VSS 0
Vprobe_517_to_VSS PROBE<517> VSS 0
Vprobe_518_to_VSS PROBE<518> VSS 0
Vprobe_519_to_VSS PROBE<519> VSS 0
Vprobe_520_to_VSS PROBE<520> VSS 0
Vprobe_521_to_VSS PROBE<521> VSS 0
Vprobe_522_to_VSS PROBE<522> VSS 0
Vprobe_523_to_VSS PROBE<523> VSS 0
Vprobe_524_to_VSS PROBE<524> VSS 0
Vprobe_525_to_VSS PROBE<525> VSS 0
Vprobe_526_to_VSS PROBE<526> VSS 0
Vprobe_527_to_VSS PROBE<527> VSS 0
Vprobe_528_to_VSS PROBE<528> VSS 0
Vprobe_529_to_VSS PROBE<529> VSS 0
Vprobe_530_to_VSS PROBE<530> VSS 0
Vprobe_533_to_VSS PROBE<533> VSS 0
Vprobe_534_to_VSS PROBE<534> VSS 0
Vprobe_535_to_VSS PROBE<535> VSS 0
Vprobe_536_to_VSS PROBE<536> VSS 0
Vprobe_537_to_VSS PROBE<537> VSS 0
Vprobe_538_to_VSS PROBE<538> VSS 0
Vprobe_539_to_VSS PROBE<539> VSS 0
Vprobe_540_to_VSS PROBE<540> VSS 0
Vprobe_541_to_VSS PROBE<541> VSS 0
Vprobe_542_to_VSS PROBE<542> VSS 0
Vprobe_543_to_VSS PROBE<543> VSS 0
Vprobe_544_to_VSS PROBE<544> VSS 0
Vprobe_545_to_VSS PROBE<545> VSS 0
Vprobe_546_to_VSS PROBE<546> VSS 0
Vprobe_547_to_VSS PROBE<547> VSS 0
Vprobe_548_to_VSS PROBE<548> VSS 0
Vprobe_549_to_VSS PROBE<549> VSS 0
Vprobe_550_to_VSS PROBE<550> VSS 0
Vprobe_551_to_VSS PROBE<551> VSS 0
Vprobe_552_to_VSS PROBE<552> VSS 0
Vprobe_553_to_VSS PROBE<553> VSS 0
Vprobe_554_to_VSS PROBE<554> VSS 0
Vprobe_555_to_VSS PROBE<555> VSS 0
Vprobe_556_to_VSS PROBE<556> VSS 0
Vprobe_557_to_VSS PROBE<557> VSS 0
Vprobe_558_to_VSS PROBE<558> VSS 0
Vprobe_559_to_VSS PROBE<559> VSS 0
Vprobe_560_to_VSS PROBE<560> VSS 0
Vprobe_561_to_VSS PROBE<561> VSS 0
Vprobe_562_to_VSS PROBE<562> VSS 0
Vprobe_563_to_VSS PROBE<563> VSS 0
Vprobe_564_to_VSS PROBE<564> VSS 0
Vprobe_565_to_VSS PROBE<565> VSS 0
Vprobe_566_to_VSS PROBE<566> VSS 0
Vprobe_567_to_VSS PROBE<567> VSS 0
Vprobe_568_to_VSS PROBE<568> VSS 0
Vprobe_569_to_VSS PROBE<569> VSS 0
Vprobe_570_to_VSS PROBE<570> VSS 0
Vprobe_571_to_VSS PROBE<571> VSS 0
Vprobe_572_to_VSS PROBE<572> VSS 0
Vprobe_573_to_VSS PROBE<573> VSS 0
Vprobe_574_to_VSS PROBE<574> VSS 0
Vprobe_575_to_VSS PROBE<575> VSS 0
Vprobe_576_to_VSS PROBE<576> VSS 0
Vprobe_577_to_VSS PROBE<577> VSS 0
Vprobe_578_to_VSS PROBE<578> VSS 0
Vprobe_579_to_VSS PROBE<579> VSS 0
Vprobe_580_to_VSS PROBE<580> VSS 0
Vprobe_581_to_VSS PROBE<581> VSS 0
Vprobe_582_to_VSS PROBE<582> VSS 0
Vprobe_583_to_VSS PROBE<583> VSS 0
Vprobe_584_to_VSS PROBE<584> VSS 0
Vprobe_585_to_VSS PROBE<585> VSS 0
Vprobe_586_to_VSS PROBE<586> VSS 0
Vprobe_587_to_VSS PROBE<587> VSS 0
Vprobe_588_to_VSS PROBE<588> VSS 0
Vprobe_589_to_VSS PROBE<589> VSS 0
Vprobe_590_to_VSS PROBE<590> VSS 0
Vprobe_591_to_VSS PROBE<591> VSS 0
Vprobe_592_to_VSS PROBE<592> VSS 0
Vprobe_593_to_VSS PROBE<593> VSS 0
Vprobe_594_to_VSS PROBE<594> VSS 0
Vprobe_595_to_VSS PROBE<595> VSS 0
Vprobe_596_to_VSS PROBE<596> VSS 0
Vprobe_597_to_VSS PROBE<597> VSS 0
Vprobe_598_to_VSS PROBE<598> VSS 0
Vprobe_599_to_VSS PROBE<599> VSS 0
Vprobe_600_to_VSS PROBE<600> VSS 0
Vprobe_601_to_VSS PROBE<601> VSS 0
Vprobe_602_to_VSS PROBE<602> VSS 0
Vprobe_603_to_VSS PROBE<603> VSS 0
Vprobe_604_to_VSS PROBE<604> VSS 0
Vprobe_605_to_VSS PROBE<605> VSS 0
Vprobe_606_to_VSS PROBE<606> VSS 0
Vprobe_607_to_VSS PROBE<607> VSS 0
Vprobe_608_to_VSS PROBE<608> VSS 0
Vprobe_609_to_VSS PROBE<609> VSS 0
Vprobe_610_to_VSS PROBE<610> VSS 0
Vprobe_611_to_VSS PROBE<611> VSS 0
Vprobe_612_to_VSS PROBE<612> VSS 0
Vprobe_613_to_VSS PROBE<613> VSS 0
Vprobe_614_to_VSS PROBE<614> VSS 0
Vprobe_615_to_VSS PROBE<615> VSS 0
Vprobe_616_to_VSS PROBE<616> VSS 0
Vprobe_617_to_VSS PROBE<617> VSS 0
Vprobe_618_to_VSS PROBE<618> VSS 0
Vprobe_619_to_VSS PROBE<619> VSS 0
Vprobe_620_to_VSS PROBE<620> VSS 0
Vprobe_621_to_VSS PROBE<621> VSS 0
Vprobe_622_to_VSS PROBE<622> VSS 0
Vprobe_623_to_VSS PROBE<623> VSS 0
Vprobe_624_to_VSS PROBE<624> VSS 0
Vprobe_625_to_VSS PROBE<625> VSS 0
Vprobe_626_to_VSS PROBE<626> VSS 0
Vprobe_627_to_VSS PROBE<627> VSS 0
Vprobe_628_to_VSS PROBE<628> VSS 0
Vprobe_629_to_VSS PROBE<629> VSS 0
Vprobe_630_to_VSS PROBE<630> VSS 0
Vprobe_631_to_VSS PROBE<631> VSS 0
Vprobe_632_to_VSS PROBE<632> VSS 0
Vprobe_633_to_VSS PROBE<633> VSS 0
Vprobe_634_to_VSS PROBE<634> VSS 0
Vprobe_635_to_VSS PROBE<635> VSS 0
Vprobe_636_to_VSS PROBE<636> VSS 0
Vprobe_637_to_VSS PROBE<637> VSS 0
Vprobe_638_to_VSS PROBE<638> VSS 0
Vprobe_639_to_VSS PROBE<639> VSS 0
Vprobe_640_to_VSS PROBE<640> VSS 0
Vprobe_641_to_VSS PROBE<641> VSS 0
Vprobe_642_to_VSS PROBE<642> VSS 0
Vprobe_643_to_VSS PROBE<643> VSS 0
Vprobe_644_to_VSS PROBE<644> VSS 0
Vprobe_645_to_VSS PROBE<645> VSS 0
Vprobe_646_to_VSS PROBE<646> VSS 0
Vprobe_647_to_VSS PROBE<647> VSS 0
Vprobe_648_to_VSS PROBE<648> VSS 0
Vprobe_649_to_VSS PROBE<649> VSS 0
Vprobe_650_to_VSS PROBE<650> VSS 0
Vprobe_651_to_VSS PROBE<651> VSS 0
Vprobe_652_to_VSS PROBE<652> VSS 0
Vprobe_653_to_VSS PROBE<653> VSS 0
Vprobe_654_to_VSS PROBE<654> VSS 0
Vprobe_655_to_VSS PROBE<655> VSS 0
Vprobe_656_to_VSS PROBE<656> VSS 0
Vprobe_657_to_VSS PROBE<657> VSS 0
Vprobe_658_to_VSS PROBE<658> VSS 0
Vprobe_659_to_VSS PROBE<659> VSS 0
Vprobe_660_to_VSS PROBE<660> VSS 0
Vprobe_661_to_VSS PROBE<661> VSS 0
Vprobe_662_to_VSS PROBE<662> VSS 0
Vprobe_663_to_VSS PROBE<663> VSS 0
Vprobe_664_to_VSS PROBE<664> VSS 0
Vprobe_665_to_VSS PROBE<665> VSS 0
Vprobe_666_to_VSS PROBE<666> VSS 0
Vprobe_667_to_VSS PROBE<667> VSS 0
Vprobe_668_to_VSS PROBE<668> VSS 0
Vprobe_669_to_VSS PROBE<669> VSS 0
Vprobe_670_to_VSS PROBE<670> VSS 0
Vprobe_671_to_VSS PROBE<671> VSS 0
Vprobe_672_to_VSS PROBE<672> VSS 0
Vprobe_673_to_VSS PROBE<673> VSS 0
Vprobe_674_to_VSS PROBE<674> VSS 0
Vprobe_675_to_VSS PROBE<675> VSS 0
Vprobe_676_to_VSS PROBE<676> VSS 0
Vprobe_677_to_VSS PROBE<677> VSS 0
Vprobe_678_to_VSS PROBE<678> VSS 0
Vprobe_679_to_VSS PROBE<679> VSS 0
Vprobe_680_to_VSS PROBE<680> VSS 0
Vprobe_681_to_VSS PROBE<681> VSS 0
Vprobe_682_to_VSS PROBE<682> VSS 0
Vprobe_683_to_VSS PROBE<683> VSS 0
Vprobe_684_to_VSS PROBE<684> VSS 0
Vprobe_685_to_VSS PROBE<685> VSS 0
Vprobe_686_to_VSS PROBE<686> VSS 0
Vprobe_687_to_VSS PROBE<687> VSS 0
Vprobe_688_to_VSS PROBE<688> VSS 0
Vprobe_689_to_VSS PROBE<689> VSS 0
Vprobe_690_to_VSS PROBE<690> VSS 0
Vprobe_691_to_VSS PROBE<691> VSS 0
Vprobe_692_to_VSS PROBE<692> VSS 0
Vprobe_693_to_VSS PROBE<693> VSS 0
Vprobe_694_to_VSS PROBE<694> VSS 0
Vprobe_695_to_VSS PROBE<695> VSS 0
Vprobe_696_to_VSS PROBE<696> VSS 0
Vprobe_697_to_VSS PROBE<697> VSS 0
Vprobe_698_to_VSS PROBE<698> VSS 0
Vprobe_699_to_VSS PROBE<699> VSS 0
Vprobe_700_to_VSS PROBE<700> VSS 0
Vprobe_701_to_VSS PROBE<701> VSS 0
Vprobe_702_to_VSS PROBE<702> VSS 0
Vprobe_703_to_VSS PROBE<703> VSS 0
Vprobe_704_to_VSS PROBE<704> VSS 0
Vprobe_705_to_VSS PROBE<705> VSS 0
Vprobe_706_to_VSS PROBE<706> VSS 0
Vprobe_707_to_VSS PROBE<707> VSS 0
Vprobe_708_to_VSS PROBE<708> VSS 0
Vprobe_709_to_VSS PROBE<709> VSS 0
Vprobe_710_to_VSS PROBE<710> VSS 0
Vprobe_711_to_VSS PROBE<711> VSS 0
Vprobe_712_to_VSS PROBE<712> VSS 0
Vprobe_713_to_VSS PROBE<713> VSS 0
Vprobe_714_to_VSS PROBE<714> VSS 0
Vprobe_715_to_VSS PROBE<715> VSS 0
Vprobe_716_to_VSS PROBE<716> VSS 0
Vprobe_717_to_VSS PROBE<717> VSS 0
Vprobe_718_to_VSS PROBE<718> VSS 0
Vprobe_719_to_VSS PROBE<719> VSS 0
Vprobe_720_to_VSS PROBE<720> VSS 0
Vprobe_721_to_VSS PROBE<721> VSS 0
Vprobe_722_to_VSS PROBE<722> VSS 0
Vprobe_723_to_VSS PROBE<723> VSS 0
Vprobe_724_to_VSS PROBE<724> VSS 0
Vprobe_725_to_VSS PROBE<725> VSS 0
Vprobe_726_to_VSS PROBE<726> VSS 0
Vprobe_727_to_VSS PROBE<727> VSS 0
Vprobe_728_to_VSS PROBE<728> VSS 0
Vprobe_729_to_VSS PROBE<729> VSS 0
Vprobe_730_to_VSS PROBE<730> VSS 0
Vprobe_731_to_VSS PROBE<731> VSS 0
Vprobe_732_to_VSS PROBE<732> VSS 0
Vprobe_733_to_VSS PROBE<733> VSS 0
Vprobe_734_to_VSS PROBE<734> VSS 0
Vprobe_735_to_VSS PROBE<735> VSS 0
Vprobe_736_to_VSS PROBE<736> VSS 0
Vprobe_737_to_VSS PROBE<737> VSS 0
Vprobe_738_to_VSS PROBE<738> VSS 0
Vprobe_739_to_VSS PROBE<739> VSS 0
Vprobe_740_to_VSS PROBE<740> VSS 0
Vprobe_741_to_VSS PROBE<741> VSS 0
Vprobe_742_to_VSS PROBE<742> VSS 0
Vprobe_743_to_VSS PROBE<743> VSS 0
Vprobe_744_to_VSS PROBE<744> VSS 0
Vprobe_745_to_VSS PROBE<745> VSS 0
Vprobe_746_to_VSS PROBE<746> VSS 0
Vprobe_747_to_VSS PROBE<747> VSS 0
Vprobe_748_to_VSS PROBE<748> VSS 0
Vprobe_749_to_VSS PROBE<749> VSS 0
Vprobe_750_to_VSS PROBE<750> VSS 0
Vprobe_751_to_VSS PROBE<751> VSS 0
Vprobe_752_to_VSS PROBE<752> VSS 0
Vprobe_753_to_VSS PROBE<753> VSS 0
Vprobe_754_to_VSS PROBE<754> VSS 0
Vprobe_755_to_VSS PROBE<755> VSS 0
Vprobe_756_to_VSS PROBE<756> VSS 0
Vprobe_757_to_VSS PROBE<757> VSS 0
Vprobe_758_to_VSS PROBE<758> VSS 0
Vprobe_759_to_VSS PROBE<759> VSS 0
Vprobe_760_to_VSS PROBE<760> VSS 0
Vprobe_761_to_VSS PROBE<761> VSS 0
Vprobe_762_to_VSS PROBE<762> VSS 0
Vprobe_763_to_VSS PROBE<763> VSS 0
Vprobe_764_to_VSS PROBE<764> VSS 0
Vprobe_765_to_VSS PROBE<765> VSS 0
Vprobe_766_to_VSS PROBE<766> VSS 0
Vprobe_767_to_VSS PROBE<767> VSS 0
Vprobe_768_to_VSS PROBE<768> VSS 0
Vprobe_769_to_VSS PROBE<769> VSS 0
Vprobe_770_to_VSS PROBE<770> VSS 0
Vprobe_771_to_VSS PROBE<771> VSS 0
Vprobe_772_to_VSS PROBE<772> VSS 0
Vprobe_773_to_VSS PROBE<773> VSS 0
Vprobe_774_to_VSS PROBE<774> VSS 0
Vprobe_775_to_VSS PROBE<775> VSS 0
Vprobe_776_to_VSS PROBE<776> VSS 0
Vprobe_777_to_VSS PROBE<777> VSS 0
Vprobe_778_to_VSS PROBE<778> VSS 0
Vprobe_779_to_VSS PROBE<779> VSS 0
Vprobe_780_to_VSS PROBE<780> VSS 0
Vprobe_781_to_VSS PROBE<781> VSS 0
Vprobe_782_to_VSS PROBE<782> VSS 0
Vprobe_783_to_VSS PROBE<783> VSS 0
Vprobe_784_to_VSS PROBE<784> VSS 0
Vprobe_785_to_VSS PROBE<785> VSS 0
Vprobe_786_to_VSS PROBE<786> VSS 0
Vprobe_787_to_VSS PROBE<787> VSS 0
Vprobe_788_to_VSS PROBE<788> VSS 0
Vprobe_789_to_VSS PROBE<789> VSS 0
Vprobe_790_to_VSS PROBE<790> VSS 0
Vprobe_792_to_VSS PROBE<792> VSS 0
Vprobe_793_to_VSS PROBE<793> VSS 0
Vprobe_794_to_VSS PROBE<794> VSS 0
Vprobe_795_to_VSS PROBE<795> VSS 0
Vprobe_796_to_VSS PROBE<796> VSS 0
Vprobe_797_to_VSS PROBE<797> VSS 0
Vprobe_798_to_VSS PROBE<798> VSS 0
Vprobe_799_to_VSS PROBE<799> VSS 0
Vprobe_800_to_VSS PROBE<800> VSS 0
Vprobe_801_to_VSS PROBE<801> VSS 0
Vprobe_802_to_VSS PROBE<802> VSS 0
Vprobe_803_to_VSS PROBE<803> VSS 0
Vprobe_804_to_VSS PROBE<804> VSS 0
Vprobe_805_to_VSS PROBE<805> VSS 0
Vprobe_806_to_VSS PROBE<806> VSS 0
Vprobe_807_to_VSS PROBE<807> VSS 0
Vprobe_808_to_VSS PROBE<808> VSS 0
Vprobe_809_to_VSS PROBE<809> VSS 0
Vprobe_810_to_VSS PROBE<810> VSS 0
Vprobe_811_to_VSS PROBE<811> VSS 0
Vprobe_812_to_VSS PROBE<812> VSS 0
Vprobe_813_to_VSS PROBE<813> VSS 0
Vprobe_814_to_VSS PROBE<814> VSS 0
Vprobe_815_to_VSS PROBE<815> VSS 0
Vprobe_817_to_VSS PROBE<817> VSS 0
Vprobe_819_to_VSS PROBE<819> VSS 0
Vprobe_820_to_VSS PROBE<820> VSS 0
Vprobe_821_to_VSS PROBE<821> VSS 0
Vprobe_822_to_VSS PROBE<822> VSS 0
Vprobe_823_to_VSS PROBE<823> VSS 0
Vprobe_824_to_VSS PROBE<824> VSS 0
Vprobe_825_to_VSS PROBE<825> VSS 0
Vprobe_826_to_VSS PROBE<826> VSS 0
Vprobe_827_to_VSS PROBE<827> VSS 0
Vprobe_828_to_VSS PROBE<828> VSS 0
Vprobe_829_to_VSS PROBE<829> VSS 0
Vprobe_830_to_VSS PROBE<830> VSS 0
Vprobe_831_to_VSS PROBE<831> VSS 0
Vprobe_832_to_VSS PROBE<832> VSS 0
Vprobe_833_to_VSS PROBE<833> VSS 0
Vprobe_834_to_VSS PROBE<834> VSS 0
Vprobe_835_to_VSS PROBE<835> VSS 0
Vprobe_836_to_VSS PROBE<836> VSS 0
Vprobe_837_to_VSS PROBE<837> VSS 0
Vprobe_838_to_VSS PROBE<838> VSS 0
Vprobe_839_to_VSS PROBE<839> VSS 0
Vprobe_840_to_VSS PROBE<840> VSS 0
Vprobe_841_to_VSS PROBE<841> VSS 0
Vprobe_842_to_VSS PROBE<842> VSS 0
Vprobe_844_to_VSS PROBE<844> VSS 0
Vprobe_846_to_VSS PROBE<846> VSS 0
Vprobe_847_to_VSS PROBE<847> VSS 0
Vprobe_848_to_VSS PROBE<848> VSS 0
Vprobe_849_to_VSS PROBE<849> VSS 0
Vprobe_850_to_VSS PROBE<850> VSS 0
Vprobe_851_to_VSS PROBE<851> VSS 0
Vprobe_852_to_VSS PROBE<852> VSS 0
Vprobe_853_to_VSS PROBE<853> VSS 0
Vprobe_854_to_VSS PROBE<854> VSS 0
Vprobe_855_to_VSS PROBE<855> VSS 0
Vprobe_856_to_VSS PROBE<856> VSS 0
Vprobe_857_to_VSS PROBE<857> VSS 0
Vprobe_858_to_VSS PROBE<858> VSS 0
Vprobe_859_to_VSS PROBE<859> VSS 0
Vprobe_860_to_VSS PROBE<860> VSS 0
Vprobe_861_to_VSS PROBE<861> VSS 0
Vprobe_862_to_VSS PROBE<862> VSS 0
Vprobe_863_to_VSS PROBE<863> VSS 0
Vprobe_864_to_VSS PROBE<864> VSS 0
Vprobe_865_to_VSS PROBE<865> VSS 0
Vprobe_866_to_VSS PROBE<866> VSS 0
Vprobe_867_to_VSS PROBE<867> VSS 0
Vprobe_868_to_VSS PROBE<868> VSS 0
Vprobe_869_to_VSS PROBE<869> VSS 0
Vprobe_871_to_VSS PROBE<871> VSS 0
Vprobe_873_to_VSS PROBE<873> VSS 0
Vprobe_874_to_VSS PROBE<874> VSS 0
Vprobe_875_to_VSS PROBE<875> VSS 0
Vprobe_876_to_VSS PROBE<876> VSS 0
Vprobe_877_to_VSS PROBE<877> VSS 0
Vprobe_878_to_VSS PROBE<878> VSS 0
Vprobe_879_to_VSS PROBE<879> VSS 0
Vprobe_880_to_VSS PROBE<880> VSS 0
Vprobe_881_to_VSS PROBE<881> VSS 0
Vprobe_882_to_VSS PROBE<882> VSS 0
Vprobe_883_to_VSS PROBE<883> VSS 0
Vprobe_884_to_VSS PROBE<884> VSS 0
Vprobe_885_to_VSS PROBE<885> VSS 0
Vprobe_886_to_VSS PROBE<886> VSS 0
Vprobe_887_to_VSS PROBE<887> VSS 0
Vprobe_888_to_VSS PROBE<888> VSS 0
Vprobe_889_to_VSS PROBE<889> VSS 0
Vprobe_890_to_VSS PROBE<890> VSS 0
Vprobe_891_to_VSS PROBE<891> VSS 0
Vprobe_892_to_VSS PROBE<892> VSS 0
Vprobe_893_to_VSS PROBE<893> VSS 0
Vprobe_894_to_VSS PROBE<894> VSS 0
Vprobe_895_to_VSS PROBE<895> VSS 0
Vprobe_896_to_VSS PROBE<896> VSS 0
Vprobe_897_to_VSS PROBE<897> VSS 0
Vprobe_898_to_VSS PROBE<898> VSS 0
Vprobe_899_to_VSS PROBE<899> VSS 0
Vprobe_900_to_VSS PROBE<900> VSS 0
Vprobe_901_to_VSS PROBE<901> VSS 0
Vprobe_902_to_VSS PROBE<902> VSS 0
Vprobe_903_to_VSS PROBE<903> VSS 0
Vprobe_904_to_VSS PROBE<904> VSS 0
Vprobe_905_to_VSS PROBE<905> VSS 0
Vprobe_906_to_VSS PROBE<906> VSS 0
Vprobe_907_to_VSS PROBE<907> VSS 0
Vprobe_908_to_VSS PROBE<908> VSS 0
Vprobe_909_to_VSS PROBE<909> VSS 0
Vprobe_910_to_VSS PROBE<910> VSS 0
Vprobe_911_to_VSS PROBE<911> VSS 0
Vprobe_912_to_VSS PROBE<912> VSS 0
Vprobe_913_to_VSS PROBE<913> VSS 0
Vprobe_914_to_VSS PROBE<914> VSS 0
Vprobe_915_to_VSS PROBE<915> VSS 0
Vprobe_916_to_VSS PROBE<916> VSS 0
Vprobe_917_to_VSS PROBE<917> VSS 0
Vprobe_918_to_VSS PROBE<918> VSS 0
Vprobe_919_to_VSS PROBE<919> VSS 0
Vprobe_920_to_VSS PROBE<920> VSS 0
Vprobe_921_to_VSS PROBE<921> VSS 0
Vprobe_922_to_VSS PROBE<922> VSS 0
Vprobe_923_to_VSS PROBE<923> VSS 0
Vprobe_924_to_VSS PROBE<924> VSS 0
Vprobe_925_to_VSS PROBE<925> VSS 0
Vprobe_927_to_VSS PROBE<927> VSS 0
Vprobe_928_to_VSS PROBE<928> VSS 0
Vprobe_929_to_VSS PROBE<929> VSS 0
Vprobe_931_to_VSS PROBE<931> VSS 0
Vprobe_933_to_VSS PROBE<933> VSS 0
Vprobe_934_to_VSS PROBE<934> VSS 0
Vprobe_935_to_VSS PROBE<935> VSS 0
Vprobe_936_to_VSS PROBE<936> VSS 0
Vprobe_937_to_VSS PROBE<937> VSS 0
Vprobe_939_to_VSS PROBE<939> VSS 0
Vprobe_941_to_VSS PROBE<941> VSS 0
Vprobe_942_to_VSS PROBE<942> VSS 0
Vprobe_943_to_VSS PROBE<943> VSS 0
Vprobe_944_to_VSS PROBE<944> VSS 0
Vprobe_945_to_VSS PROBE<945> VSS 0
Vprobe_946_to_VSS PROBE<946> VSS 0
Vprobe_947_to_VSS PROBE<947> VSS 0
Vprobe_948_to_VSS PROBE<948> VSS 0
Vprobe_949_to_VSS PROBE<949> VSS 0
Vprobe_950_to_VSS PROBE<950> VSS 0
Vprobe_951_to_VSS PROBE<951> VSS 0
Vprobe_952_to_VSS PROBE<952> VSS 0
Vprobe_953_to_VSS PROBE<953> VSS 0
Vprobe_954_to_VSS PROBE<954> VSS 0
Vprobe_955_to_VSS PROBE<955> VSS 0
Vprobe_956_to_VSS PROBE<956> VSS 0
Vprobe_957_to_VSS PROBE<957> VSS 0
Vprobe_958_to_VSS PROBE<958> VSS 0
Vprobe_959_to_VSS PROBE<959> VSS 0
Vprobe_960_to_VSS PROBE<960> VSS 0
Vprobe_961_to_VSS PROBE<961> VSS 0
Vprobe_962_to_VSS PROBE<962> VSS 0
Vprobe_963_to_VSS PROBE<963> VSS 0
Vprobe_964_to_VSS PROBE<964> VSS 0
Vprobe_965_to_VSS PROBE<965> VSS 0
Vprobe_966_to_VSS PROBE<966> VSS 0
Vprobe_967_to_VSS PROBE<967> VSS 0
Vprobe_968_to_VSS PROBE<968> VSS 0
Vprobe_969_to_VSS PROBE<969> VSS 0
Vprobe_970_to_VSS PROBE<970> VSS 0
Vprobe_971_to_VSS PROBE<971> VSS 0
Vprobe_972_to_VSS PROBE<972> VSS 0
Vprobe_973_to_VSS PROBE<973> VSS 0
Vprobe_974_to_VSS PROBE<974> VSS 0
Vprobe_975_to_VSS PROBE<975> VSS 0
Vprobe_976_to_VSS PROBE<976> VSS 0
Vprobe_977_to_VSS PROBE<977> VSS 0
Vprobe_978_to_VSS PROBE<978> VSS 0
Vprobe_979_to_VSS PROBE<979> VSS 0
Vprobe_980_to_VSS PROBE<980> VSS 0
Vprobe_981_to_VSS PROBE<981> VSS 0
Vprobe_982_to_VSS PROBE<982> VSS 0
Vprobe_983_to_VSS PROBE<983> VSS 0
Vprobe_984_to_VSS PROBE<984> VSS 0
Vprobe_985_to_VSS PROBE<985> VSS 0
Vprobe_986_to_VSS PROBE<986> VSS 0
Vprobe_987_to_VSS PROBE<987> VSS 0
Vprobe_988_to_VSS PROBE<988> VSS 0
Vprobe_989_to_VSS PROBE<989> VSS 0
Vprobe_990_to_VSS PROBE<990> VSS 0
Vprobe_991_to_VSS PROBE<991> VSS 0
Vprobe_992_to_VSS PROBE<992> VSS 0
Vprobe_993_to_VSS PROBE<993> VSS 0
Vprobe_994_to_VSS PROBE<994> VSS 0
Vprobe_995_to_VSS PROBE<995> VSS 0
Vprobe_996_to_VSS PROBE<996> VSS 0
Vprobe_997_to_VSS PROBE<997> VSS 0
Vprobe_998_to_VSS PROBE<998> VSS 0
Vprobe_999_to_VSS PROBE<999> VSS 0
Vprobe_1000_to_VSS PROBE<1000> VSS 0
Vprobe_1001_to_VSS PROBE<1001> VSS 0
Vprobe_1002_to_VSS PROBE<1002> VSS 0
Vprobe_1003_to_VSS PROBE<1003> VSS 0
Vprobe_1004_to_VSS PROBE<1004> VSS 0
Vprobe_1005_to_VSS PROBE<1005> VSS 0
Vprobe_1006_to_VSS PROBE<1006> VSS 0
Vprobe_1007_to_VSS PROBE<1007> VSS 0
Vprobe_1008_to_VSS PROBE<1008> VSS 0
Vprobe_1009_to_VSS PROBE<1009> VSS 0
Vprobe_1010_to_VSS PROBE<1010> VSS 0
Vprobe_1011_to_VSS PROBE<1011> VSS 0
Vprobe_1012_to_VSS PROBE<1012> VSS 0
Vprobe_1013_to_VSS PROBE<1013> VSS 0
Vprobe_1014_to_VSS PROBE<1014> VSS 0
Vprobe_1015_to_VSS PROBE<1015> VSS 0
Vprobe_1016_to_VSS PROBE<1016> VSS 0
Vprobe_1017_to_VSS PROBE<1017> VSS 0
Vprobe_1018_to_VSS PROBE<1018> VSS 0
Vprobe_1019_to_VSS PROBE<1019> VSS 0
Vprobe_1020_to_VSS PROBE<1020> VSS 0
Vprobe_1021_to_VSS PROBE<1021> VSS 0
Vprobe_1022_to_VSS PROBE<1022> VSS 0
Vprobe_1023_to_VSS PROBE<1023> VSS 0
Vprobe_1024_to_VSS PROBE<1024> VSS 0
Vprobe_1025_to_VSS PROBE<1025> VSS 0
Vprobe_1026_to_VSS PROBE<1026> VSS 0
Vprobe_1027_to_VSS PROBE<1027> VSS 0
Vprobe_1028_to_VSS PROBE<1028> VSS 0
Vprobe_1029_to_VSS PROBE<1029> VSS 0
Vprobe_1030_to_VSS PROBE<1030> VSS 0
Vprobe_1031_to_VSS PROBE<1031> VSS 0
Vprobe_1032_to_VSS PROBE<1032> VSS 0
Vprobe_1033_to_VSS PROBE<1033> VSS 0
Vprobe_1034_to_VSS PROBE<1034> VSS 0
Vprobe_1035_to_VSS PROBE<1035> VSS 0
Vprobe_1036_to_VSS PROBE<1036> VSS 0
Vprobe_1037_to_VSS PROBE<1037> VSS 0
Vprobe_1038_to_VSS PROBE<1038> VSS 0
Vprobe_1039_to_VSS PROBE<1039> VSS 0
Vprobe_1040_to_VSS PROBE<1040> VSS 0
Vprobe_1041_to_VSS PROBE<1041> VSS 0
Vprobe_1042_to_VSS PROBE<1042> VSS 0
Vprobe_1043_to_VSS PROBE<1043> VSS 0
Vprobe_1044_to_VSS PROBE<1044> VSS 0
Vprobe_1045_to_VSS PROBE<1045> VSS 0
Vprobe_1046_to_VSS PROBE<1046> VSS 0
Vprobe_1047_to_VSS PROBE<1047> VSS 0
Vprobe_1048_to_VSS PROBE<1048> VSS 0
Vprobe_1049_to_VSS PROBE<1049> VSS 0
Vprobe_1050_to_VSS PROBE<1050> VSS 0
Vprobe_1051_to_VSS PROBE<1051> VSS 0
Vprobe_1052_to_VSS PROBE<1052> VSS 0
Vprobe_1053_to_VSS PROBE<1053> VSS 0
Vprobe_1054_to_VSS PROBE<1054> VSS 0
Vprobe_1055_to_VSS PROBE<1055> VSS 0
Vprobe_1056_to_VSS PROBE<1056> VSS 0
Vprobe_1057_to_VSS PROBE<1057> VSS 0
Vprobe_1058_to_VSS PROBE<1058> VSS 0
Vprobe_1059_to_VSS PROBE<1059> VSS 0
Vprobe_1060_to_VSS PROBE<1060> VSS 0
Vprobe_1061_to_VSS PROBE<1061> VSS 0
Vprobe_1062_to_VSS PROBE<1062> VSS 0
Vprobe_1063_to_VSS PROBE<1063> VSS 0
Vprobe_1064_to_VSS PROBE<1064> VSS 0
Vprobe_1065_to_VSS PROBE<1065> VSS 0
Vprobe_1066_to_VSS PROBE<1066> VSS 0
Vprobe_1067_to_VSS PROBE<1067> VSS 0
Vprobe_1068_to_VSS PROBE<1068> VSS 0
Vprobe_1069_to_VSS PROBE<1069> VSS 0
Vprobe_1070_to_VSS PROBE<1070> VSS 0
Vprobe_1071_to_VSS PROBE<1071> VSS 0
Vprobe_1072_to_VSS PROBE<1072> VSS 0
Vprobe_1073_to_VSS PROBE<1073> VSS 0
Vprobe_1074_to_VSS PROBE<1074> VSS 0
Vprobe_1075_to_VSS PROBE<1075> VSS 0
Vprobe_1076_to_VSS PROBE<1076> VSS 0
Vprobe_1077_to_VSS PROBE<1077> VSS 0
Vprobe_1078_to_VSS PROBE<1078> VSS 0
Vprobe_1079_to_VSS PROBE<1079> VSS 0
Vprobe_1080_to_VSS PROBE<1080> VSS 0
Vprobe_1081_to_VSS PROBE<1081> VSS 0
Vprobe_1082_to_VSS PROBE<1082> VSS 0
Vprobe_1083_to_VSS PROBE<1083> VSS 0
Vprobe_1084_to_VSS PROBE<1084> VSS 0
Vprobe_1085_to_VSS PROBE<1085> VSS 0
Vprobe_1086_to_VSS PROBE<1086> VSS 0
Vprobe_1087_to_VSS PROBE<1087> VSS 0
Vprobe_1088_to_VSS PROBE<1088> VSS 0
Vprobe_1089_to_VSS PROBE<1089> VSS 0
Vprobe_1090_to_VSS PROBE<1090> VSS 0
Vprobe_1091_to_VSS PROBE<1091> VSS 0
Vprobe_1092_to_VSS PROBE<1092> VSS 0
Vprobe_1093_to_VSS PROBE<1093> VSS 0
Vprobe_1094_to_VSS PROBE<1094> VSS 0
Vprobe_1095_to_VSS PROBE<1095> VSS 0
Vprobe_1096_to_VSS PROBE<1096> VSS 0
Vprobe_1097_to_VSS PROBE<1097> VSS 0
Vprobe_1098_to_VSS PROBE<1098> VSS 0
Vprobe_1099_to_VSS PROBE<1099> VSS 0
Vprobe_1100_to_VSS PROBE<1100> VSS 0
Vprobe_1101_to_VSS PROBE<1101> VSS 0
Vprobe_1102_to_VSS PROBE<1102> VSS 0
Vprobe_1103_to_VSS PROBE<1103> VSS 0
Vprobe_1104_to_VSS PROBE<1104> VSS 0
Vprobe_1105_to_VSS PROBE<1105> VSS 0
Vprobe_1106_to_VSS PROBE<1106> VSS 0
Vprobe_1107_to_VSS PROBE<1107> VSS 0
Vprobe_1108_to_VSS PROBE<1108> VSS 0
Vprobe_1109_to_VSS PROBE<1109> VSS 0
Vprobe_1110_to_VSS PROBE<1110> VSS 0
Vprobe_1111_to_VSS PROBE<1111> VSS 0
Vprobe_1112_to_VSS PROBE<1112> VSS 0
Vprobe_1113_to_VSS PROBE<1113> VSS 0
Vprobe_1114_to_VSS PROBE<1114> VSS 0
Vprobe_1115_to_VSS PROBE<1115> VSS 0
Vprobe_1116_to_VSS PROBE<1116> VSS 0
Vprobe_1117_to_VSS PROBE<1117> VSS 0
Vprobe_1118_to_VSS PROBE<1118> VSS 0
Vprobe_1119_to_VSS PROBE<1119> VSS 0
Vprobe_1120_to_VSS PROBE<1120> VSS 0
Vprobe_1121_to_VSS PROBE<1121> VSS 0
Vprobe_1122_to_VSS PROBE<1122> VSS 0
Vprobe_1123_to_VSS PROBE<1123> VSS 0
Vprobe_1124_to_VSS PROBE<1124> VSS 0
Vprobe_1125_to_VSS PROBE<1125> VSS 0
Vprobe_1126_to_VSS PROBE<1126> VSS 0
Vprobe_1127_to_VSS PROBE<1127> VSS 0
Vprobe_1128_to_VSS PROBE<1128> VSS 0
Vprobe_1129_to_VSS PROBE<1129> VSS 0
Vprobe_1130_to_VSS PROBE<1130> VSS 0
Vprobe_1131_to_VSS PROBE<1131> VSS 0
Vprobe_1132_to_VSS PROBE<1132> VSS 0
Vprobe_1133_to_VSS PROBE<1133> VSS 0
Vprobe_1134_to_VSS PROBE<1134> VSS 0
Vprobe_1135_to_VSS PROBE<1135> VSS 0
Vprobe_1136_to_VSS PROBE<1136> VSS 0
Vprobe_1137_to_VSS PROBE<1137> VSS 0
Vprobe_1138_to_VSS PROBE<1138> VSS 0
Vprobe_1139_to_VSS PROBE<1139> VSS 0
Vprobe_1140_to_VSS PROBE<1140> VSS 0
Vprobe_1141_to_VSS PROBE<1141> VSS 0
Vprobe_1142_to_VSS PROBE<1142> VSS 0
Vprobe_1143_to_VSS PROBE<1143> VSS 0
Vprobe_1144_to_VSS PROBE<1144> VSS 0
Vprobe_1145_to_VSS PROBE<1145> VSS 0
Vprobe_1146_to_VSS PROBE<1146> VSS 0
Vprobe_1147_to_VSS PROBE<1147> VSS 0
Vprobe_1148_to_VSS PROBE<1148> VSS 0
Vprobe_1149_to_VSS PROBE<1149> VSS 0
Vprobe_1150_to_VSS PROBE<1150> VSS 0
Vprobe_1151_to_VSS PROBE<1151> VSS 0
Vprobe_1152_to_VSS PROBE<1152> VSS 0
Vprobe_1153_to_VSS PROBE<1153> VSS 0
Vprobe_1154_to_VSS PROBE<1154> VSS 0
Vprobe_1155_to_VSS PROBE<1155> VSS 0
Vprobe_1156_to_VSS PROBE<1156> VSS 0
Vprobe_1157_to_VSS PROBE<1157> VSS 0
Vprobe_1158_to_VSS PROBE<1158> VSS 0
Vprobe_1159_to_VSS PROBE<1159> VSS 0
Vprobe_1160_to_VSS PROBE<1160> VSS 0
Vprobe_1161_to_VSS PROBE<1161> VSS 0
Vprobe_1162_to_VSS PROBE<1162> VSS 0
Vprobe_1163_to_VSS PROBE<1163> VSS 0
Vprobe_1164_to_VSS PROBE<1164> VSS 0
Vprobe_1165_to_VSS PROBE<1165> VSS 0
Vprobe_1166_to_VSS PROBE<1166> VSS 0
Vprobe_1167_to_VSS PROBE<1167> VSS 0
Vprobe_1168_to_VSS PROBE<1168> VSS 0
Vprobe_1169_to_VSS PROBE<1169> VSS 0
Vprobe_1170_to_VSS PROBE<1170> VSS 0
Vprobe_1171_to_VSS PROBE<1171> VSS 0
Vprobe_1172_to_VSS PROBE<1172> VSS 0
Vprobe_1173_to_VSS PROBE<1173> VSS 0
Vprobe_1174_to_VSS PROBE<1174> VSS 0
Vprobe_1175_to_VSS PROBE<1175> VSS 0
Vprobe_1176_to_VSS PROBE<1176> VSS 0
Vprobe_1177_to_VSS PROBE<1177> VSS 0
Vprobe_1178_to_VSS PROBE<1178> VSS 0
Vprobe_1179_to_VSS PROBE<1179> VSS 0
Vprobe_1180_to_VSS PROBE<1180> VSS 0
Vprobe_1181_to_VSS PROBE<1181> VSS 0
Vprobe_1182_to_VSS PROBE<1182> VSS 0
Vprobe_1183_to_VSS PROBE<1183> VSS 0
Vprobe_1184_to_VSS PROBE<1184> VSS 0
Vprobe_1185_to_VSS PROBE<1185> VSS 0
Vprobe_1186_to_VSS PROBE<1186> VSS 0
Vprobe_1187_to_VSS PROBE<1187> VSS 0
Vprobe_1188_to_VSS PROBE<1188> VSS 0
Vprobe_1189_to_VSS PROBE<1189> VSS 0
Vprobe_1190_to_VSS PROBE<1190> VSS 0
Vprobe_1191_to_VSS PROBE<1191> VSS 0
Vprobe_1192_to_VSS PROBE<1192> VSS 0
Vprobe_1193_to_VSS PROBE<1193> VSS 0
Vprobe_1194_to_VSS PROBE<1194> VSS 0
Vprobe_1195_to_VSS PROBE<1195> VSS 0
Vprobe_1196_to_VSS PROBE<1196> VSS 0
Vprobe_1197_to_VSS PROBE<1197> VSS 0
Vprobe_1198_to_VSS PROBE<1198> VSS 0
Vprobe_1199_to_VSS PROBE<1199> VSS 0
Vprobe_1200_to_VSS PROBE<1200> VSS 0
Vprobe_1203_to_VSS PROBE<1203> VSS 0
Vprobe_1204_to_VSS PROBE<1204> VSS 0
Vprobe_1205_to_VSS PROBE<1205> VSS 0
Vprobe_1206_to_VSS PROBE<1206> VSS 0
Vprobe_1207_to_VSS PROBE<1207> VSS 0
Vprobe_1208_to_VSS PROBE<1208> VSS 0
Vprobe_1209_to_VSS PROBE<1209> VSS 0
Vprobe_1210_to_VSS PROBE<1210> VSS 0
Vprobe_1211_to_VSS PROBE<1211> VSS 0
Vprobe_1212_to_VSS PROBE<1212> VSS 0
Vprobe_1213_to_VSS PROBE<1213> VSS 0
Vprobe_1214_to_VSS PROBE<1214> VSS 0
Vprobe_1215_to_VSS PROBE<1215> VSS 0
Vprobe_1216_to_VSS PROBE<1216> VSS 0
Vprobe_1217_to_VSS PROBE<1217> VSS 0
Vprobe_1218_to_VSS PROBE<1218> VSS 0
Vprobe_1219_to_VSS PROBE<1219> VSS 0
Vprobe_1220_to_VSS PROBE<1220> VSS 0
Vprobe_1221_to_VSS PROBE<1221> VSS 0
Vprobe_1222_to_VSS PROBE<1222> VSS 0
Vprobe_1223_to_VSS PROBE<1223> VSS 0
Vprobe_1224_to_VSS PROBE<1224> VSS 0
Vprobe_1225_to_VSS PROBE<1225> VSS 0
Vprobe_1226_to_VSS PROBE<1226> VSS 0
Vprobe_1227_to_VSS PROBE<1227> VSS 0
Vprobe_1228_to_VSS PROBE<1228> VSS 0
Vprobe_1229_to_VSS PROBE<1229> VSS 0
Vprobe_1230_to_VSS PROBE<1230> VSS 0
Vprobe_1231_to_VSS PROBE<1231> VSS 0
Vprobe_1232_to_VSS PROBE<1232> VSS 0
Vprobe_1233_to_VSS PROBE<1233> VSS 0
Vprobe_1234_to_VSS PROBE<1234> VSS 0
Vprobe_1235_to_VSS PROBE<1235> VSS 0
Vprobe_1236_to_VSS PROBE<1236> VSS 0
Vprobe_1237_to_VSS PROBE<1237> VSS 0
Vprobe_1238_to_VSS PROBE<1238> VSS 0
Vprobe_1239_to_VSS PROBE<1239> VSS 0
Vprobe_1240_to_VSS PROBE<1240> VSS 0
Vprobe_1241_to_VSS PROBE<1241> VSS 0
Vprobe_1242_to_VSS PROBE<1242> VSS 0
Vprobe_1244_to_VSS PROBE<1244> VSS 0
Vprobe_1246_to_VSS PROBE<1246> VSS 0
Vprobe_1247_to_VSS PROBE<1247> VSS 0
Vprobe_1248_to_VSS PROBE<1248> VSS 0
Vprobe_1249_to_VSS PROBE<1249> VSS 0
Vprobe_1250_to_VSS PROBE<1250> VSS 0
Vprobe_1251_to_VSS PROBE<1251> VSS 0
Vprobe_1252_to_VSS PROBE<1252> VSS 0
Vprobe_1253_to_VSS PROBE<1253> VSS 0
Vprobe_1254_to_VSS PROBE<1254> VSS 0
Vprobe_1255_to_VSS PROBE<1255> VSS 0
Vprobe_1256_to_VSS PROBE<1256> VSS 0
Vprobe_1257_to_VSS PROBE<1257> VSS 0
Vprobe_1258_to_VSS PROBE<1258> VSS 0
Vprobe_1259_to_VSS PROBE<1259> VSS 0
Vprobe_1260_to_VSS PROBE<1260> VSS 0
Vprobe_1261_to_VSS PROBE<1261> VSS 0
Vprobe_1262_to_VSS PROBE<1262> VSS 0
Vprobe_1263_to_VSS PROBE<1263> VSS 0
Vprobe_1264_to_VSS PROBE<1264> VSS 0
Vprobe_1265_to_VSS PROBE<1265> VSS 0
Vprobe_1266_to_VSS PROBE<1266> VSS 0
Vprobe_1267_to_VSS PROBE<1267> VSS 0
Vprobe_1268_to_VSS PROBE<1268> VSS 0
Vprobe_1269_to_VSS PROBE<1269> VSS 0
Vprobe_1271_to_VSS PROBE<1271> VSS 0
Vprobe_1272_to_VSS PROBE<1272> VSS 0
Vprobe_1274_to_VSS PROBE<1274> VSS 0
Vprobe_1275_to_VSS PROBE<1275> VSS 0
Vprobe_1276_to_VSS PROBE<1276> VSS 0
Vprobe_1277_to_VSS PROBE<1277> VSS 0
Vprobe_1278_to_VSS PROBE<1278> VSS 0
Vprobe_1279_to_VSS PROBE<1279> VSS 0
Vprobe_1280_to_VSS PROBE<1280> VSS 0
Vprobe_1281_to_VSS PROBE<1281> VSS 0
Vprobe_1282_to_VSS PROBE<1282> VSS 0
Vprobe_1283_to_VSS PROBE<1283> VSS 0
Vprobe_1284_to_VSS PROBE<1284> VSS 0
Vprobe_1285_to_VSS PROBE<1285> VSS 0
Vprobe_1286_to_VSS PROBE<1286> VSS 0
Vprobe_1287_to_VSS PROBE<1287> VSS 0
Vprobe_1288_to_VSS PROBE<1288> VSS 0
Vprobe_1289_to_VSS PROBE<1289> VSS 0
Vprobe_1290_to_VSS PROBE<1290> VSS 0
Vprobe_1291_to_VSS PROBE<1291> VSS 0
Vprobe_1292_to_VSS PROBE<1292> VSS 0
Vprobe_1293_to_VSS PROBE<1293> VSS 0
Vprobe_1294_to_VSS PROBE<1294> VSS 0
Vprobe_1295_to_VSS PROBE<1295> VSS 0
Vprobe_1296_to_VSS PROBE<1296> VSS 0
Vprobe_1297_to_VSS PROBE<1297> VSS 0
Vprobe_1299_to_VSS PROBE<1299> VSS 0
Vprobe_1301_to_VSS PROBE<1301> VSS 0
Vprobe_1302_to_VSS PROBE<1302> VSS 0
Vprobe_1304_to_VSS PROBE<1304> VSS 0
Vprobe_1305_to_VSS PROBE<1305> VSS 0
Vprobe_1306_to_VSS PROBE<1306> VSS 0
Vprobe_1307_to_VSS PROBE<1307> VSS 0
Vprobe_1308_to_VSS PROBE<1308> VSS 0
Vprobe_1309_to_VSS PROBE<1309> VSS 0
Vprobe_1310_to_VSS PROBE<1310> VSS 0
Vprobe_1311_to_VSS PROBE<1311> VSS 0
Vprobe_1312_to_VSS PROBE<1312> VSS 0
Vprobe_1313_to_VSS PROBE<1313> VSS 0
Vprobe_1314_to_VSS PROBE<1314> VSS 0
Vprobe_1315_to_VSS PROBE<1315> VSS 0
Vprobe_1316_to_VSS PROBE<1316> VSS 0
Vprobe_1317_to_VSS PROBE<1317> VSS 0
Vprobe_1318_to_VSS PROBE<1318> VSS 0
Vprobe_1319_to_VSS PROBE<1319> VSS 0
Vprobe_1320_to_VSS PROBE<1320> VSS 0
Vprobe_1321_to_VSS PROBE<1321> VSS 0
Vprobe_1322_to_VSS PROBE<1322> VSS 0
Vprobe_1323_to_VSS PROBE<1323> VSS 0
Vprobe_1324_to_VSS PROBE<1324> VSS 0
Vprobe_1325_to_VSS PROBE<1325> VSS 0
Vprobe_1326_to_VSS PROBE<1326> VSS 0
Vprobe_1327_to_VSS PROBE<1327> VSS 0
Vprobe_1329_to_VSS PROBE<1329> VSS 0
Vprobe_1331_to_VSS PROBE<1331> VSS 0
Vprobe_1332_to_VSS PROBE<1332> VSS 0
Vprobe_1333_to_VSS PROBE<1333> VSS 0
Vprobe_1334_to_VSS PROBE<1334> VSS 0
Vprobe_1335_to_VSS PROBE<1335> VSS 0
Vprobe_1336_to_VSS PROBE<1336> VSS 0
Vprobe_1337_to_VSS PROBE<1337> VSS 0
Vprobe_1338_to_VSS PROBE<1338> VSS 0
Vprobe_1339_to_VSS PROBE<1339> VSS 0
Vprobe_1340_to_VSS PROBE<1340> VSS 0
Vprobe_1341_to_VSS PROBE<1341> VSS 0
Vprobe_1342_to_VSS PROBE<1342> VSS 0
Vprobe_1343_to_VSS PROBE<1343> VSS 0
Vprobe_1344_to_VSS PROBE<1344> VSS 0
Vprobe_1345_to_VSS PROBE<1345> VSS 0
Vprobe_1346_to_VSS PROBE<1346> VSS 0
Vprobe_1347_to_VSS PROBE<1347> VSS 0
Vprobe_1348_to_VSS PROBE<1348> VSS 0
Vprobe_1349_to_VSS PROBE<1349> VSS 0
Vprobe_1350_to_VSS PROBE<1350> VSS 0
Vprobe_1351_to_VSS PROBE<1351> VSS 0
Vprobe_1352_to_VSS PROBE<1352> VSS 0
Vprobe_1353_to_VSS PROBE<1353> VSS 0
Vprobe_1354_to_VSS PROBE<1354> VSS 0
Vprobe_1355_to_VSS PROBE<1355> VSS 0
Vprobe_1356_to_VSS PROBE<1356> VSS 0
Vprobe_1357_to_VSS PROBE<1357> VSS 0
Vprobe_1358_to_VSS PROBE<1358> VSS 0
Vprobe_1359_to_VSS PROBE<1359> VSS 0
Vprobe_1360_to_VSS PROBE<1360> VSS 0
Vprobe_1361_to_VSS PROBE<1361> VSS 0
Vprobe_1362_to_VSS PROBE<1362> VSS 0
Vprobe_1363_to_VSS PROBE<1363> VSS 0
Vprobe_1364_to_VSS PROBE<1364> VSS 0
Vprobe_1365_to_VSS PROBE<1365> VSS 0
Vprobe_1366_to_VSS PROBE<1366> VSS 0
Vprobe_1367_to_VSS PROBE<1367> VSS 0
Vprobe_1368_to_VSS PROBE<1368> VSS 0
Vprobe_1369_to_VSS PROBE<1369> VSS 0
Vprobe_1370_to_VSS PROBE<1370> VSS 0
Vprobe_1372_to_VSS PROBE<1372> VSS 0
Vprobe_1374_to_VSS PROBE<1374> VSS 0
Vprobe_1375_to_VSS PROBE<1375> VSS 0
Vprobe_1376_to_VSS PROBE<1376> VSS 0
Vprobe_1377_to_VSS PROBE<1377> VSS 0
Vprobe_1378_to_VSS PROBE<1378> VSS 0
Vprobe_1379_to_VSS PROBE<1379> VSS 0
Vprobe_1380_to_VSS PROBE<1380> VSS 0
Vprobe_1381_to_VSS PROBE<1381> VSS 0
Vprobe_1382_to_VSS PROBE<1382> VSS 0
Vprobe_1383_to_VSS PROBE<1383> VSS 0
Vprobe_1384_to_VSS PROBE<1384> VSS 0
Vprobe_1385_to_VSS PROBE<1385> VSS 0
Vprobe_1386_to_VSS PROBE<1386> VSS 0
Vprobe_1388_to_VSS PROBE<1388> VSS 0
Vprobe_1390_to_VSS PROBE<1390> VSS 0
Vprobe_1391_to_VSS PROBE<1391> VSS 0
Vprobe_1392_to_VSS PROBE<1392> VSS 0
Vprobe_1393_to_VSS PROBE<1393> VSS 0
Vprobe_1394_to_VSS PROBE<1394> VSS 0
Vprobe_1395_to_VSS PROBE<1395> VSS 0
Vprobe_1396_to_VSS PROBE<1396> VSS 0
Vprobe_1397_to_VSS PROBE<1397> VSS 0
Vprobe_1398_to_VSS PROBE<1398> VSS 0
Vprobe_1399_to_VSS PROBE<1399> VSS 0
Vprobe_1400_to_VSS PROBE<1400> VSS 0
Vprobe_1401_to_VSS PROBE<1401> VSS 0
Vprobe_1402_to_VSS PROBE<1402> VSS 0
Vprobe_1404_to_VSS PROBE<1404> VSS 0
Vprobe_1406_to_VSS PROBE<1406> VSS 0
Vprobe_1407_to_VSS PROBE<1407> VSS 0
Vprobe_1408_to_VSS PROBE<1408> VSS 0
Vprobe_1409_to_VSS PROBE<1409> VSS 0
Vprobe_1410_to_VSS PROBE<1410> VSS 0
Vprobe_1411_to_VSS PROBE<1411> VSS 0
Vprobe_1412_to_VSS PROBE<1412> VSS 0
Vprobe_1413_to_VSS PROBE<1413> VSS 0
Vprobe_1414_to_VSS PROBE<1414> VSS 0
Vprobe_1415_to_VSS PROBE<1415> VSS 0
Vprobe_1416_to_VSS PROBE<1416> VSS 0
Vprobe_1417_to_VSS PROBE<1417> VSS 0
Vprobe_1418_to_VSS PROBE<1418> VSS 0
Vprobe_1419_to_VSS PROBE<1419> VSS 0
Vprobe_1420_to_VSS PROBE<1420> VSS 0
Vprobe_1421_to_VSS PROBE<1421> VSS 0
Vprobe_1422_to_VSS PROBE<1422> VSS 0
Vprobe_1423_to_VSS PROBE<1423> VSS 0
Vprobe_1424_to_VSS PROBE<1424> VSS 0
Vprobe_1425_to_VSS PROBE<1425> VSS 0
Vprobe_1426_to_VSS PROBE<1426> VSS 0
Vprobe_1429_to_VSS PROBE<1429> VSS 0
Vprobe_1430_to_VSS PROBE<1430> VSS 0
Vprobe_1431_to_VSS PROBE<1431> VSS 0
Vprobe_1432_to_VSS PROBE<1432> VSS 0
Vprobe_1433_to_VSS PROBE<1433> VSS 0
Vprobe_1434_to_VSS PROBE<1434> VSS 0
Vprobe_1435_to_VSS PROBE<1435> VSS 0
Vprobe_1436_to_VSS PROBE<1436> VSS 0
Vprobe_1437_to_VSS PROBE<1437> VSS 0
Vprobe_1438_to_VSS PROBE<1438> VSS 0
Vprobe_1439_to_VSS PROBE<1439> VSS 0
Vprobe_1440_to_VSS PROBE<1440> VSS 0
Vprobe_1441_to_VSS PROBE<1441> VSS 0
Vprobe_1442_to_VSS PROBE<1442> VSS 0
Vprobe_1443_to_VSS PROBE<1443> VSS 0
Vprobe_1444_to_VSS PROBE<1444> VSS 0
Vprobe_1445_to_VSS PROBE<1445> VSS 0
Vprobe_1446_to_VSS PROBE<1446> VSS 0
Vprobe_1447_to_VSS PROBE<1447> VSS 0
Vprobe_1448_to_VSS PROBE<1448> VSS 0
Vprobe_1449_to_VSS PROBE<1449> VSS 0
Vprobe_1450_to_VSS PROBE<1450> VSS 0
Vprobe_1451_to_VSS PROBE<1451> VSS 0
Vprobe_1452_to_VSS PROBE<1452> VSS 0
Vprobe_1453_to_VSS PROBE<1453> VSS 0
Vprobe_1454_to_VSS PROBE<1454> VSS 0
Vprobe_1455_to_VSS PROBE<1455> VSS 0
Vprobe_1456_to_VSS PROBE<1456> VSS 0
Vprobe_1457_to_VSS PROBE<1457> VSS 0
Vprobe_1458_to_VSS PROBE<1458> VSS 0
Vprobe_1459_to_VSS PROBE<1459> VSS 0
Vprobe_1460_to_VSS PROBE<1460> VSS 0
Vprobe_1461_to_VSS PROBE<1461> VSS 0
Vprobe_1462_to_VSS PROBE<1462> VSS 0
Vprobe_1463_to_VSS PROBE<1463> VSS 0
Vprobe_1464_to_VSS PROBE<1464> VSS 0
Vprobe_1465_to_VSS PROBE<1465> VSS 0
Vprobe_1466_to_VSS PROBE<1466> VSS 0
Vprobe_1467_to_VSS PROBE<1467> VSS 0
Vprobe_1468_to_VSS PROBE<1468> VSS 0
Vprobe_1469_to_VSS PROBE<1469> VSS 0
Vprobe_1470_to_VSS PROBE<1470> VSS 0
Vprobe_1471_to_VSS PROBE<1471> VSS 0
Vprobe_1472_to_VSS PROBE<1472> VSS 0
Vprobe_1473_to_VSS PROBE<1473> VSS 0
Vprobe_1474_to_VSS PROBE<1474> VSS 0
Vprobe_1475_to_VSS PROBE<1475> VSS 0
Vprobe_1476_to_VSS PROBE<1476> VSS 0
Vprobe_1477_to_VSS PROBE<1477> VSS 0
Vprobe_1478_to_VSS PROBE<1478> VSS 0
Vprobe_1481_to_VSS PROBE<1481> VSS 0
Vprobe_1482_to_VSS PROBE<1482> VSS 0
Vprobe_1483_to_VSS PROBE<1483> VSS 0
Vprobe_1484_to_VSS PROBE<1484> VSS 0
Vprobe_1485_to_VSS PROBE<1485> VSS 0
Vprobe_1486_to_VSS PROBE<1486> VSS 0
Vprobe_1487_to_VSS PROBE<1487> VSS 0
Vprobe_1488_to_VSS PROBE<1488> VSS 0
Vprobe_1489_to_VSS PROBE<1489> VSS 0
Vprobe_1490_to_VSS PROBE<1490> VSS 0
Vprobe_1491_to_VSS PROBE<1491> VSS 0
Vprobe_1492_to_VSS PROBE<1492> VSS 0
Vprobe_1493_to_VSS PROBE<1493> VSS 0
Vprobe_1494_to_VSS PROBE<1494> VSS 0
Vprobe_1495_to_VSS PROBE<1495> VSS 0
Vprobe_1496_to_VSS PROBE<1496> VSS 0
Vprobe_1497_to_VSS PROBE<1497> VSS 0
Vprobe_1498_to_VSS PROBE<1498> VSS 0
Vprobe_1499_to_VSS PROBE<1499> VSS 0
Vprobe_1500_to_VSS PROBE<1500> VSS 0
Vprobe_1501_to_VSS PROBE<1501> VSS 0
Vprobe_1502_to_VSS PROBE<1502> VSS 0
Vprobe_1503_to_VSS PROBE<1503> VSS 0
Vprobe_1504_to_VSS PROBE<1504> VSS 0
Vprobe_1505_to_VSS PROBE<1505> VSS 0
Vprobe_1506_to_VSS PROBE<1506> VSS 0
Vprobe_1507_to_VSS PROBE<1507> VSS 0
Vprobe_1508_to_VSS PROBE<1508> VSS 0
Vprobe_1509_to_VSS PROBE<1509> VSS 0
Vprobe_1510_to_VSS PROBE<1510> VSS 0
Vprobe_1511_to_VSS PROBE<1511> VSS 0
Vprobe_1512_to_VSS PROBE<1512> VSS 0
Vprobe_1513_to_VSS PROBE<1513> VSS 0
Vprobe_1514_to_VSS PROBE<1514> VSS 0
Vprobe_1515_to_VSS PROBE<1515> VSS 0
Vprobe_1516_to_VSS PROBE<1516> VSS 0
Vprobe_1517_to_VSS PROBE<1517> VSS 0
Vprobe_1518_to_VSS PROBE<1518> VSS 0
Vprobe_1519_to_VSS PROBE<1519> VSS 0
Vprobe_1520_to_VSS PROBE<1520> VSS 0
Vprobe_1521_to_VSS PROBE<1521> VSS 0
Vprobe_1522_to_VSS PROBE<1522> VSS 0
Vprobe_1523_to_VSS PROBE<1523> VSS 0
Vprobe_1524_to_VSS PROBE<1524> VSS 0
Vprobe_1525_to_VSS PROBE<1525> VSS 0
Vprobe_1526_to_VSS PROBE<1526> VSS 0
Vprobe_1527_to_VSS PROBE<1527> VSS 0
Vprobe_1528_to_VSS PROBE<1528> VSS 0
Vprobe_1529_to_VSS PROBE<1529> VSS 0
Vprobe_1530_to_VSS PROBE<1530> VSS 0
Vprobe_1531_to_VSS PROBE<1531> VSS 0
Vprobe_1532_to_VSS PROBE<1532> VSS 0
Vprobe_1533_to_VSS PROBE<1533> VSS 0
Vprobe_1534_to_VSS PROBE<1534> VSS 0
Vprobe_1535_to_VSS PROBE<1535> VSS 0
Vprobe_1536_to_VSS PROBE<1536> VSS 0
Vprobe_1537_to_VSS PROBE<1537> VSS 0
Vprobe_1538_to_VSS PROBE<1538> VSS 0
Vprobe_1539_to_VSS PROBE<1539> VSS 0
Vprobe_1540_to_VSS PROBE<1540> VSS 0
Vprobe_1541_to_VSS PROBE<1541> VSS 0
Vprobe_1542_to_VSS PROBE<1542> VSS 0
Vprobe_1543_to_VSS PROBE<1543> VSS 0
Vprobe_1544_to_VSS PROBE<1544> VSS 0
Vprobe_1545_to_VSS PROBE<1545> VSS 0
Vprobe_1546_to_VSS PROBE<1546> VSS 0
Vprobe_1547_to_VSS PROBE<1547> VSS 0
Vprobe_1548_to_VSS PROBE<1548> VSS 0
Vprobe_1549_to_VSS PROBE<1549> VSS 0
Vprobe_1550_to_VSS PROBE<1550> VSS 0
Vprobe_1551_to_VSS PROBE<1551> VSS 0
Vprobe_1552_to_VSS PROBE<1552> VSS 0
Vprobe_1553_to_VSS PROBE<1553> VSS 0
Vprobe_1554_to_VSS PROBE<1554> VSS 0
Vprobe_1555_to_VSS PROBE<1555> VSS 0
Vprobe_1556_to_VSS PROBE<1556> VSS 0
Vprobe_1557_to_VSS PROBE<1557> VSS 0
Vprobe_1558_to_VSS PROBE<1558> VSS 0
Vprobe_1559_to_VSS PROBE<1559> VSS 0
Vprobe_1560_to_VSS PROBE<1560> VSS 0
Vprobe_1561_to_VSS PROBE<1561> VSS 0
Vprobe_1562_to_VSS PROBE<1562> VSS 0
Vprobe_1563_to_VSS PROBE<1563> VSS 0
Vprobe_1564_to_VSS PROBE<1564> VSS 0
Vprobe_1565_to_VSS PROBE<1565> VSS 0
Vprobe_1566_to_VSS PROBE<1566> VSS 0
Vprobe_1567_to_VSS PROBE<1567> VSS 0
Vprobe_1568_to_VSS PROBE<1568> VSS 0
Vprobe_1569_to_VSS PROBE<1569> VSS 0
Vprobe_1570_to_VSS PROBE<1570> VSS 0
Vprobe_1571_to_VSS PROBE<1571> VSS 0
Vprobe_1572_to_VSS PROBE<1572> VSS 0
Vprobe_1573_to_VSS PROBE<1573> VSS 0
Vprobe_1574_to_VSS PROBE<1574> VSS 0
Vprobe_1575_to_VSS PROBE<1575> VSS 0
Vprobe_1576_to_VSS PROBE<1576> VSS 0
Vprobe_1577_to_VSS PROBE<1577> VSS 0
Vprobe_1578_to_VSS PROBE<1578> VSS 0
Vprobe_1579_to_VSS PROBE<1579> VSS 0
Vprobe_1580_to_VSS PROBE<1580> VSS 0
Vprobe_1581_to_VSS PROBE<1581> VSS 0
Vprobe_1582_to_VSS PROBE<1582> VSS 0
Vprobe_1583_to_VSS PROBE<1583> VSS 0
Vprobe_1584_to_VSS PROBE<1584> VSS 0
Vprobe_1585_to_VSS PROBE<1585> VSS 0
Vprobe_1586_to_VSS PROBE<1586> VSS 0
Vprobe_1587_to_VSS PROBE<1587> VSS 0
Vprobe_1588_to_VSS PROBE<1588> VSS 0
Vprobe_1589_to_VSS PROBE<1589> VSS 0
Vprobe_1590_to_VSS PROBE<1590> VSS 0
Vprobe_1591_to_VSS PROBE<1591> VSS 0
Vprobe_1592_to_VSS PROBE<1592> VSS 0
Vprobe_1593_to_VSS PROBE<1593> VSS 0
Vprobe_1594_to_VSS PROBE<1594> VSS 0
Vprobe_1595_to_VSS PROBE<1595> VSS 0
Vprobe_1596_to_VSS PROBE<1596> VSS 0
Vprobe_1597_to_VSS PROBE<1597> VSS 0
Vprobe_1598_to_VSS PROBE<1598> VSS 0
Vprobe_1599_to_VSS PROBE<1599> VSS 0
Vprobe_1600_to_VSS PROBE<1600> VSS 0
Vprobe_1601_to_VSS PROBE<1601> VSS 0
Vprobe_1602_to_VSS PROBE<1602> VSS 0
Vprobe_1603_to_VSS PROBE<1603> VSS 0
Vprobe_1604_to_VSS PROBE<1604> VSS 0
Vprobe_1605_to_VSS PROBE<1605> VSS 0
Vprobe_1606_to_VSS PROBE<1606> VSS 0
Vprobe_1607_to_VSS PROBE<1607> VSS 0
Vprobe_1608_to_VSS PROBE<1608> VSS 0
Vprobe_1609_to_VSS PROBE<1609> VSS 0
Vprobe_1610_to_VSS PROBE<1610> VSS 0
Vprobe_1611_to_VSS PROBE<1611> VSS 0
Vprobe_1612_to_VSS PROBE<1612> VSS 0
Vprobe_1613_to_VSS PROBE<1613> VSS 0
Vprobe_1614_to_VSS PROBE<1614> VSS 0
Vprobe_1615_to_VSS PROBE<1615> VSS 0
Vprobe_1616_to_VSS PROBE<1616> VSS 0
Vprobe_1617_to_VSS PROBE<1617> VSS 0
Vprobe_1618_to_VSS PROBE<1618> VSS 0
Vprobe_1619_to_VSS PROBE<1619> VSS 0
Vprobe_1620_to_VSS PROBE<1620> VSS 0
Vprobe_1621_to_VSS PROBE<1621> VSS 0
Vprobe_1622_to_VSS PROBE<1622> VSS 0
Vprobe_1623_to_VSS PROBE<1623> VSS 0
Vprobe_1624_to_VSS PROBE<1624> VSS 0
Vprobe_1625_to_VSS PROBE<1625> VSS 0
Vprobe_1626_to_VSS PROBE<1626> VSS 0
Vprobe_1627_to_VSS PROBE<1627> VSS 0
Vprobe_1628_to_VSS PROBE<1628> VSS 0
Vprobe_1629_to_VSS PROBE<1629> VSS 0
Vprobe_1630_to_VSS PROBE<1630> VSS 0
Vprobe_1631_to_VSS PROBE<1631> VSS 0
Vprobe_1632_to_VSS PROBE<1632> VSS 0
Vprobe_1633_to_VSS PROBE<1633> VSS 0
Vprobe_1634_to_VSS PROBE<1634> VSS 0
Vprobe_1635_to_VSS PROBE<1635> VSS 0
Vprobe_1636_to_VSS PROBE<1636> VSS 0
Vprobe_1637_to_VSS PROBE<1637> VSS 0
Vprobe_1638_to_VSS PROBE<1638> VSS 0
Vprobe_1639_to_VSS PROBE<1639> VSS 0
Vprobe_1640_to_VSS PROBE<1640> VSS 0
Vprobe_1641_to_VSS PROBE<1641> VSS 0
Vprobe_1642_to_VSS PROBE<1642> VSS 0
Vprobe_1643_to_VSS PROBE<1643> VSS 0
Vprobe_1644_to_VSS PROBE<1644> VSS 0
Vprobe_1645_to_VSS PROBE<1645> VSS 0
Vprobe_1646_to_VSS PROBE<1646> VSS 0
Vprobe_1647_to_VSS PROBE<1647> VSS 0
Vprobe_1648_to_VSS PROBE<1648> VSS 0
Vprobe_1649_to_VSS PROBE<1649> VSS 0
Vprobe_1650_to_VSS PROBE<1650> VSS 0
Vprobe_1651_to_VSS PROBE<1651> VSS 0
Vprobe_1652_to_VSS PROBE<1652> VSS 0
Vprobe_1653_to_VSS PROBE<1653> VSS 0
Vprobe_1654_to_VSS PROBE<1654> VSS 0
Vprobe_1655_to_VSS PROBE<1655> VSS 0
Vprobe_1656_to_VSS PROBE<1656> VSS 0
Vprobe_1657_to_VSS PROBE<1657> VSS 0
Vprobe_1658_to_VSS PROBE<1658> VSS 0
Vprobe_1659_to_VSS PROBE<1659> VSS 0
Vprobe_1660_to_VSS PROBE<1660> VSS 0
Vprobe_1661_to_VSS PROBE<1661> VSS 0
Vprobe_1662_to_VSS PROBE<1662> VSS 0
Vprobe_1663_to_VSS PROBE<1663> VSS 0
Vprobe_1664_to_VSS PROBE<1664> VSS 0
Vprobe_1665_to_VSS PROBE<1665> VSS 0
Vprobe_1666_to_VSS PROBE<1666> VSS 0
Vprobe_1667_to_VSS PROBE<1667> VSS 0
Vprobe_1668_to_VSS PROBE<1668> VSS 0
Vprobe_1669_to_VSS PROBE<1669> VSS 0
Vprobe_1670_to_VSS PROBE<1670> VSS 0
Vprobe_1671_to_VSS PROBE<1671> VSS 0
Vprobe_1672_to_VSS PROBE<1672> VSS 0
Vprobe_1673_to_VSS PROBE<1673> VSS 0
Vprobe_1674_to_VSS PROBE<1674> VSS 0
Vprobe_1675_to_VSS PROBE<1675> VSS 0
Vprobe_1676_to_VSS PROBE<1676> VSS 0
Vprobe_1677_to_VSS PROBE<1677> VSS 0
Vprobe_1678_to_VSS PROBE<1678> VSS 0
Vprobe_1679_to_VSS PROBE<1679> VSS 0
Vprobe_1680_to_VSS PROBE<1680> VSS 0
Vprobe_1681_to_VSS PROBE<1681> VSS 0
Vprobe_1682_to_VSS PROBE<1682> VSS 0
Vprobe_1683_to_VSS PROBE<1683> VSS 0
Vprobe_1684_to_VSS PROBE<1684> VSS 0
Vprobe_1685_to_VSS PROBE<1685> VSS 0
Vprobe_1686_to_VSS PROBE<1686> VSS 0
Vprobe_1687_to_VSS PROBE<1687> VSS 0
Vprobe_1688_to_VSS PROBE<1688> VSS 0
Vprobe_1689_to_VSS PROBE<1689> VSS 0
Vprobe_1690_to_VSS PROBE<1690> VSS 0
Vprobe_1693_to_VSS PROBE<1693> VSS 0
Vprobe_1694_to_VSS PROBE<1694> VSS 0
Vprobe_1695_to_VSS PROBE<1695> VSS 0
Vprobe_1696_to_VSS PROBE<1696> VSS 0
Vprobe_1697_to_VSS PROBE<1697> VSS 0
Vprobe_1698_to_VSS PROBE<1698> VSS 0
Vprobe_1699_to_VSS PROBE<1699> VSS 0
Vprobe_1700_to_VSS PROBE<1700> VSS 0
Vprobe_1701_to_VSS PROBE<1701> VSS 0
Vprobe_1702_to_VSS PROBE<1702> VSS 0
Vprobe_1703_to_VSS PROBE<1703> VSS 0
Vprobe_1704_to_VSS PROBE<1704> VSS 0
Vprobe_1705_to_VSS PROBE<1705> VSS 0
Vprobe_1706_to_VSS PROBE<1706> VSS 0
Vprobe_1707_to_VSS PROBE<1707> VSS 0
Vprobe_1708_to_VSS PROBE<1708> VSS 0
Vprobe_1709_to_VSS PROBE<1709> VSS 0
Vprobe_1710_to_VSS PROBE<1710> VSS 0
Vprobe_1711_to_VSS PROBE<1711> VSS 0
Vprobe_1712_to_VSS PROBE<1712> VSS 0
Vprobe_1713_to_VSS PROBE<1713> VSS 0
Vprobe_1714_to_VSS PROBE<1714> VSS 0
Vprobe_1715_to_VSS PROBE<1715> VSS 0
Vprobe_1716_to_VSS PROBE<1716> VSS 0
Vprobe_1717_to_VSS PROBE<1717> VSS 0
Vprobe_1718_to_VSS PROBE<1718> VSS 0
Vprobe_1719_to_VSS PROBE<1719> VSS 0
Vprobe_1720_to_VSS PROBE<1720> VSS 0
Vprobe_1721_to_VSS PROBE<1721> VSS 0
Vprobe_1722_to_VSS PROBE<1722> VSS 0
Vprobe_1723_to_VSS PROBE<1723> VSS 0
Vprobe_1725_to_VSS PROBE<1725> VSS 0
Vprobe_1726_to_VSS PROBE<1726> VSS 0
Vprobe_1727_to_VSS PROBE<1727> VSS 0
Vprobe_1728_to_VSS PROBE<1728> VSS 0
Vprobe_1729_to_VSS PROBE<1729> VSS 0
Vprobe_1730_to_VSS PROBE<1730> VSS 0
Vprobe_1731_to_VSS PROBE<1731> VSS 0
Vprobe_1732_to_VSS PROBE<1732> VSS 0
Vprobe_1733_to_VSS PROBE<1733> VSS 0
Vprobe_1734_to_VSS PROBE<1734> VSS 0
Vprobe_1735_to_VSS PROBE<1735> VSS 0
Vprobe_1736_to_VSS PROBE<1736> VSS 0
Vprobe_1737_to_VSS PROBE<1737> VSS 0
Vprobe_1738_to_VSS PROBE<1738> VSS 0
Vprobe_1739_to_VSS PROBE<1739> VSS 0
Vprobe_1740_to_VSS PROBE<1740> VSS 0
Vprobe_1741_to_VSS PROBE<1741> VSS 0
Vprobe_1742_to_VSS PROBE<1742> VSS 0
Vprobe_1743_to_VSS PROBE<1743> VSS 0
Vprobe_1744_to_VSS PROBE<1744> VSS 0
Vprobe_1745_to_VSS PROBE<1745> VSS 0
Vprobe_1746_to_VSS PROBE<1746> VSS 0
Vprobe_1747_to_VSS PROBE<1747> VSS 0
Vprobe_1748_to_VSS PROBE<1748> VSS 0
Vprobe_1749_to_VSS PROBE<1749> VSS 0
Vprobe_1750_to_VSS PROBE<1750> VSS 0
Vprobe_1751_to_VSS PROBE<1751> VSS 0
Vprobe_1752_to_VSS PROBE<1752> VSS 0
Vprobe_1753_to_VSS PROBE<1753> VSS 0
Vprobe_1754_to_VSS PROBE<1754> VSS 0
Vprobe_1755_to_VSS PROBE<1755> VSS 0
Vprobe_1756_to_VSS PROBE<1756> VSS 0
Vprobe_1757_to_VSS PROBE<1757> VSS 0
Vprobe_1758_to_VSS PROBE<1758> VSS 0
Vprobe_1759_to_VSS PROBE<1759> VSS 0
Vprobe_1760_to_VSS PROBE<1760> VSS 0
Vprobe_1761_to_VSS PROBE<1761> VSS 0
Vprobe_1762_to_VSS PROBE<1762> VSS 0
Vprobe_1763_to_VSS PROBE<1763> VSS 0
Vprobe_1764_to_VSS PROBE<1764> VSS 0
Vprobe_1765_to_VSS PROBE<1765> VSS 0
Vprobe_1766_to_VSS PROBE<1766> VSS 0
Vprobe_1767_to_VSS PROBE<1767> VSS 0
Vprobe_1768_to_VSS PROBE<1768> VSS 0
Vprobe_1769_to_VSS PROBE<1769> VSS 0
Vprobe_1770_to_VSS PROBE<1770> VSS 0
Vprobe_1771_to_VSS PROBE<1771> VSS 0
Vprobe_1772_to_VSS PROBE<1772> VSS 0
Vprobe_1773_to_VSS PROBE<1773> VSS 0
Vprobe_1775_to_VSS PROBE<1775> VSS 0
Vprobe_1776_to_VSS PROBE<1776> VSS 0
Vprobe_1777_to_VSS PROBE<1777> VSS 0
Vprobe_1778_to_VSS PROBE<1778> VSS 0
Vprobe_1779_to_VSS PROBE<1779> VSS 0
Vprobe_1780_to_VSS PROBE<1780> VSS 0
Vprobe_1781_to_VSS PROBE<1781> VSS 0
Vprobe_1782_to_VSS PROBE<1782> VSS 0
Vprobe_1783_to_VSS PROBE<1783> VSS 0
Vprobe_1784_to_VSS PROBE<1784> VSS 0
Vprobe_1785_to_VSS PROBE<1785> VSS 0
Vprobe_1786_to_VSS PROBE<1786> VSS 0
Vprobe_1787_to_VSS PROBE<1787> VSS 0
Vprobe_1788_to_VSS PROBE<1788> VSS 0
Vprobe_1789_to_VSS PROBE<1789> VSS 0
Vprobe_1790_to_VSS PROBE<1790> VSS 0
Vprobe_1791_to_VSS PROBE<1791> VSS 0
Vprobe_1792_to_VSS PROBE<1792> VSS 0
Vprobe_1793_to_VSS PROBE<1793> VSS 0
Vprobe_1794_to_VSS PROBE<1794> VSS 0
Vprobe_1795_to_VSS PROBE<1795> VSS 0
Vprobe_1796_to_VSS PROBE<1796> VSS 0
Vprobe_1797_to_VSS PROBE<1797> VSS 0
Vprobe_1798_to_VSS PROBE<1798> VSS 0
Vprobe_1799_to_VSS PROBE<1799> VSS 0
Vprobe_1800_to_VSS PROBE<1800> VSS 0
Vprobe_1801_to_VSS PROBE<1801> VSS 0
Vprobe_1802_to_VSS PROBE<1802> VSS 0
Vprobe_1803_to_VSS PROBE<1803> VSS 0
Vprobe_1804_to_VSS PROBE<1804> VSS 0
Vprobe_1805_to_VSS PROBE<1805> VSS 0
Vprobe_1806_to_VSS PROBE<1806> VSS 0
Vprobe_1807_to_VSS PROBE<1807> VSS 0
Vprobe_1808_to_VSS PROBE<1808> VSS 0
Vprobe_1809_to_VSS PROBE<1809> VSS 0
Vprobe_1810_to_VSS PROBE<1810> VSS 0
Vprobe_1811_to_VSS PROBE<1811> VSS 0
Vprobe_1812_to_VSS PROBE<1812> VSS 0
Vprobe_1813_to_VSS PROBE<1813> VSS 0
Vprobe_1814_to_VSS PROBE<1814> VSS 0
Vprobe_1815_to_VSS PROBE<1815> VSS 0
Vprobe_1816_to_VSS PROBE<1816> VSS 0
Vprobe_1817_to_VSS PROBE<1817> VSS 0
Vprobe_1818_to_VSS PROBE<1818> VSS 0
Vprobe_1819_to_VSS PROBE<1819> VSS 0
Vprobe_1820_to_VSS PROBE<1820> VSS 0
Vprobe_1821_to_VSS PROBE<1821> VSS 0
Vprobe_1822_to_VSS PROBE<1822> VSS 0
Vprobe_1823_to_VSS PROBE<1823> VSS 0
Vprobe_1824_to_VSS PROBE<1824> VSS 0
Vprobe_1825_to_VSS PROBE<1825> VSS 0
Vprobe_1826_to_VSS PROBE<1826> VSS 0
Vprobe_1827_to_VSS PROBE<1827> VSS 0
Vprobe_1828_to_VSS PROBE<1828> VSS 0
Vprobe_1829_to_VSS PROBE<1829> VSS 0
Vprobe_1830_to_VSS PROBE<1830> VSS 0
Vprobe_1831_to_VSS PROBE<1831> VSS 0
Vprobe_1832_to_VSS PROBE<1832> VSS 0
Vprobe_1833_to_VSS PROBE<1833> VSS 0
Vprobe_1834_to_VSS PROBE<1834> VSS 0
Vprobe_1835_to_VSS PROBE<1835> VSS 0
Vprobe_1836_to_VSS PROBE<1836> VSS 0
Vprobe_1837_to_VSS PROBE<1837> VSS 0
Vprobe_1838_to_VSS PROBE<1838> VSS 0
Vprobe_1839_to_VSS PROBE<1839> VSS 0
Vprobe_1840_to_VSS PROBE<1840> VSS 0
Vprobe_1841_to_VSS PROBE<1841> VSS 0
Vprobe_1842_to_VSS PROBE<1842> VSS 0
Vprobe_1843_to_VSS PROBE<1843> VSS 0
Vprobe_1844_to_VSS PROBE<1844> VSS 0
Vprobe_1845_to_VSS PROBE<1845> VSS 0
Vprobe_1846_to_VSS PROBE<1846> VSS 0
Vprobe_1848_to_VSS PROBE<1848> VSS 0
Vprobe_1849_to_VSS PROBE<1849> VSS 0
Vprobe_1850_to_VSS PROBE<1850> VSS 0
Vprobe_1851_to_VSS PROBE<1851> VSS 0
Vprobe_1853_to_VSS PROBE<1853> VSS 0
Vprobe_1855_to_VSS PROBE<1855> VSS 0
Vprobe_1856_to_VSS PROBE<1856> VSS 0
Vprobe_1857_to_VSS PROBE<1857> VSS 0
Vprobe_1858_to_VSS PROBE<1858> VSS 0
Vprobe_1860_to_VSS PROBE<1860> VSS 0
Vprobe_1862_to_VSS PROBE<1862> VSS 0
Vprobe_1863_to_VSS PROBE<1863> VSS 0
Vprobe_1864_to_VSS PROBE<1864> VSS 0
Vprobe_1866_to_VSS PROBE<1866> VSS 0
Vprobe_1867_to_VSS PROBE<1867> VSS 0
Vprobe_1868_to_VSS PROBE<1868> VSS 0
Vprobe_1869_to_VSS PROBE<1869> VSS 0
Vprobe_1870_to_VSS PROBE<1870> VSS 0
Vprobe_1871_to_VSS PROBE<1871> VSS 0
Vprobe_1872_to_VSS PROBE<1872> VSS 0
Vprobe_1873_to_VSS PROBE<1873> VSS 0
Vprobe_1874_to_VSS PROBE<1874> VSS 0
Vprobe_1875_to_VSS PROBE<1875> VSS 0
Vprobe_1876_to_VSS PROBE<1876> VSS 0
Vprobe_1877_to_VSS PROBE<1877> VSS 0
Vprobe_1878_to_VSS PROBE<1878> VSS 0
Vprobe_1879_to_VSS PROBE<1879> VSS 0
Vprobe_1880_to_VSS PROBE<1880> VSS 0
Vprobe_1881_to_VSS PROBE<1881> VSS 0
Vprobe_1882_to_VSS PROBE<1882> VSS 0
Vprobe_1883_to_VSS PROBE<1883> VSS 0
Vprobe_1884_to_VSS PROBE<1884> VSS 0
Vprobe_1885_to_VSS PROBE<1885> VSS 0
Vprobe_1886_to_VSS PROBE<1886> VSS 0
Vprobe_1888_to_VSS PROBE<1888> VSS 0
.ENDS
