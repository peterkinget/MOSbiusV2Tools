*

simulator lang=spice

* Generated PK_set_sizes netlist 
*   for ../../examples/all_transistors_4x_sizes.json 
*   on 2025-05-06 18:22:54

.SUBCKT PK_set_sizes_2 PROBE<1889> PROBE<1890> PROBE<1891> PROBE<1892> PROBE<1893>
+  PROBE<1894> PROBE<1895> PROBE<1896> PROBE<1897> PROBE<1898> PROBE<1899>
+  PROBE<1900> PROBE<1901> PROBE<1902> PROBE<1903> PROBE<1904> PROBE<1905>
+  PROBE<1906> PROBE<1907> PROBE<1908> PROBE<1909> PROBE<1910> PROBE<1911>
+  PROBE<1912> PROBE<1913> PROBE<1914> PROBE<1915> PROBE<1916> PROBE<1917>
+  PROBE<1918> PROBE<1919> PROBE<1920> PROBE<1921> PROBE<1922> PROBE<1923>
+  PROBE<1924> PROBE<1925> PROBE<1926> PROBE<1927> PROBE<1928> PROBE<1929>
+  PROBE<1930> PROBE<1931> PROBE<1932> PROBE<1933> PROBE<1934> PROBE<1935>
+  PROBE<1936> PROBE<1937> PROBE<1938> PROBE<1939> PROBE<1940> PROBE<1941>
+  PROBE<1942> PROBE<1943> PROBE<1944> PROBE<1945> PROBE<1946> PROBE<1947>
+  PROBE<1948> PROBE<1949> PROBE<1950> PROBE<1951> PROBE<1952> PROBE<1953>
+  PROBE<1954> PROBE<1955> PROBE<1956> PROBE<1957> PROBE<1958> PROBE<1959>
+  PROBE<1960> PROBE<1961> PROBE<1962> PROBE<1963> PROBE<1964> PROBE<1965>
+  PROBE<1966> PROBE<1967> PROBE<1968> PROBE<1969> PROBE<1970> PROBE<1971>
+  PROBE<1972> PROBE<1973> PROBE<1974> PROBE<1975> PROBE<1976> PROBE<1977>
+  PROBE<1978> PROBE<1979> PROBE<1980> PROBE<1981> PROBE<1982> PROBE<1983>
+  PROBE<1984> PROBE<1985> PROBE<1986> PROBE<1987> PROBE<1988> PROBE<1989>
+  PROBE<1990> PROBE<1991> PROBE<1992> PROBE<1993> PROBE<1994> PROBE<1995>
+  PROBE<1996> PROBE<1997> PROBE<1998> PROBE<1999> PROBE<2000> PROBE<2001>
+  PROBE<2002> PROBE<2003> PROBE<2004> PROBE<2005> PROBE<2006> PROBE<2007>
+  PROBE<2008> VDD VSS

* Device: CC_N Size: 4 
V_CC_N_1934 PROBE<1934> VSS 0
V_CC_N_1935 PROBE<1935> VSS 0
V_CC_N_1936 PROBE<1936> VDD 0
V_CC_N_1937 PROBE<1937> VSS 0
V_CC_N_1938 PROBE<1938> VSS 0

* Device: CC_P Size: 4 
V_CC_P_1994 PROBE<1994> VSS 0
V_CC_P_1995 PROBE<1995> VSS 0
V_CC_P_1996 PROBE<1996> VDD 0
V_CC_P_1997 PROBE<1997> VSS 0
V_CC_P_1998 PROBE<1998> VSS 0

* Device: DCC1_N_L Size: 4 
V_DCC1_N_L_1914 PROBE<1914> VSS 0
V_DCC1_N_L_1915 PROBE<1915> VSS 0
V_DCC1_N_L_1916 PROBE<1916> VDD 0
V_DCC1_N_L_1917 PROBE<1917> VSS 0
V_DCC1_N_L_1918 PROBE<1918> VSS 0

* Device: DCC1_N_R Size: 4 
V_DCC1_N_R_1919 PROBE<1919> VSS 0
V_DCC1_N_R_1920 PROBE<1920> VSS 0
V_DCC1_N_R_1921 PROBE<1921> VDD 0
V_DCC1_N_R_1922 PROBE<1922> VSS 0
V_DCC1_N_R_1923 PROBE<1923> VSS 0

* Device: DCC1_P_L Size: 4 
V_DCC1_P_L_1889 PROBE<1889> VSS 0
V_DCC1_P_L_1890 PROBE<1890> VSS 0
V_DCC1_P_L_1891 PROBE<1891> VDD 0
V_DCC1_P_L_1892 PROBE<1892> VSS 0
V_DCC1_P_L_1893 PROBE<1893> VSS 0

* Device: DCC1_P_R Size: 4 
V_DCC1_P_R_1894 PROBE<1894> VSS 0
V_DCC1_P_R_1895 PROBE<1895> VSS 0
V_DCC1_P_R_1896 PROBE<1896> VDD 0
V_DCC1_P_R_1897 PROBE<1897> VSS 0
V_DCC1_P_R_1898 PROBE<1898> VSS 0

* Device: DCC2_N_L Size: 4 
V_DCC2_N_L_1939 PROBE<1939> VSS 0
V_DCC2_N_L_1940 PROBE<1940> VSS 0
V_DCC2_N_L_1941 PROBE<1941> VDD 0
V_DCC2_N_L_1942 PROBE<1942> VSS 0
V_DCC2_N_L_1943 PROBE<1943> VSS 0

* Device: DCC2_N_R Size: 4 
V_DCC2_N_R_1944 PROBE<1944> VSS 0
V_DCC2_N_R_1945 PROBE<1945> VSS 0
V_DCC2_N_R_1946 PROBE<1946> VDD 0
V_DCC2_N_R_1947 PROBE<1947> VSS 0
V_DCC2_N_R_1948 PROBE<1948> VSS 0

* Device: DCC2_P_L Size: 4 
V_DCC2_P_L_1904 PROBE<1904> VSS 0
V_DCC2_P_L_1905 PROBE<1905> VSS 0
V_DCC2_P_L_1906 PROBE<1906> VDD 0
V_DCC2_P_L_1907 PROBE<1907> VSS 0
V_DCC2_P_L_1908 PROBE<1908> VSS 0

* Device: DCC2_P_R Size: 4 
V_DCC2_P_R_1909 PROBE<1909> VSS 0
V_DCC2_P_R_1910 PROBE<1910> VSS 0
V_DCC2_P_R_1911 PROBE<1911> VDD 0
V_DCC2_P_R_1912 PROBE<1912> VSS 0
V_DCC2_P_R_1913 PROBE<1913> VSS 0

* Device: DCC3_N_L Size: 4 
V_DCC3_N_L_1949 PROBE<1949> VSS 0
V_DCC3_N_L_1950 PROBE<1950> VSS 0
V_DCC3_N_L_1951 PROBE<1951> VDD 0
V_DCC3_N_L_1952 PROBE<1952> VSS 0
V_DCC3_N_L_1953 PROBE<1953> VSS 0

* Device: DCC3_N_R Size: 4 
V_DCC3_N_R_1954 PROBE<1954> VSS 0
V_DCC3_N_R_1955 PROBE<1955> VSS 0
V_DCC3_N_R_1956 PROBE<1956> VDD 0
V_DCC3_N_R_1957 PROBE<1957> VSS 0
V_DCC3_N_R_1958 PROBE<1958> VSS 0

* Device: DCC3_P_L Size: 4 
V_DCC3_P_L_1924 PROBE<1924> VSS 0
V_DCC3_P_L_1925 PROBE<1925> VSS 0
V_DCC3_P_L_1926 PROBE<1926> VDD 0
V_DCC3_P_L_1927 PROBE<1927> VSS 0
V_DCC3_P_L_1928 PROBE<1928> VSS 0

* Device: DCC3_P_R Size: 4 
V_DCC3_P_R_1929 PROBE<1929> VSS 0
V_DCC3_P_R_1930 PROBE<1930> VSS 0
V_DCC3_P_R_1931 PROBE<1931> VDD 0
V_DCC3_P_R_1932 PROBE<1932> VSS 0
V_DCC3_P_R_1933 PROBE<1933> VSS 0

* Device: DCC4_N_L Size: 4 
V_DCC4_N_L_1999 PROBE<1999> VSS 0
V_DCC4_N_L_2000 PROBE<2000> VSS 0
V_DCC4_N_L_2001 PROBE<2001> VDD 0
V_DCC4_N_L_2002 PROBE<2002> VSS 0
V_DCC4_N_L_2003 PROBE<2003> VSS 0

* Device: DCC4_N_R Size: 4 
V_DCC4_N_R_2004 PROBE<2004> VSS 0
V_DCC4_N_R_2005 PROBE<2005> VSS 0
V_DCC4_N_R_2006 PROBE<2006> VDD 0
V_DCC4_N_R_2007 PROBE<2007> VSS 0
V_DCC4_N_R_2008 PROBE<2008> VSS 0

* Device: DCC4_P_L Size: 4 
V_DCC4_P_L_1964 PROBE<1964> VSS 0
V_DCC4_P_L_1965 PROBE<1965> VSS 0
V_DCC4_P_L_1966 PROBE<1966> VDD 0
V_DCC4_P_L_1967 PROBE<1967> VSS 0
V_DCC4_P_L_1968 PROBE<1968> VSS 0

* Device: DCC4_P_R Size: 4 
V_DCC4_P_R_1969 PROBE<1969> VSS 0
V_DCC4_P_R_1970 PROBE<1970> VSS 0
V_DCC4_P_R_1971 PROBE<1971> VDD 0
V_DCC4_P_R_1972 PROBE<1972> VSS 0
V_DCC4_P_R_1973 PROBE<1973> VSS 0

* Device: DINV1_L Size: 4 
V_DINV1_L_1974 PROBE<1974> VSS 0
V_DINV1_L_1975 PROBE<1975> VSS 0
V_DINV1_L_1976 PROBE<1976> VDD 0
V_DINV1_L_1977 PROBE<1977> VSS 0
V_DINV1_L_1978 PROBE<1978> VSS 0

* Device: DINV1_R Size: 4 
V_DINV1_R_1979 PROBE<1979> VSS 0
V_DINV1_R_1980 PROBE<1980> VSS 0
V_DINV1_R_1981 PROBE<1981> VDD 0
V_DINV1_R_1982 PROBE<1982> VSS 0
V_DINV1_R_1983 PROBE<1983> VSS 0

* Device: DINV2_L Size: 4 
V_DINV2_L_1984 PROBE<1984> VSS 0
V_DINV2_L_1985 PROBE<1985> VSS 0
V_DINV2_L_1986 PROBE<1986> VDD 0
V_DINV2_L_1987 PROBE<1987> VSS 0
V_DINV2_L_1988 PROBE<1988> VSS 0

* Device: DINV2_R Size: 4 
V_DINV2_R_1989 PROBE<1989> VSS 0
V_DINV2_R_1990 PROBE<1990> VSS 0
V_DINV2_R_1991 PROBE<1991> VDD 0
V_DINV2_R_1992 PROBE<1992> VSS 0
V_DINV2_R_1993 PROBE<1993> VSS 0

* Device: OTA_N Size: 4 
V_OTA_N_1899 PROBE<1899> VSS 0
V_OTA_N_1900 PROBE<1900> VSS 0
V_OTA_N_1901 PROBE<1901> VDD 0
V_OTA_N_1902 PROBE<1902> VSS 0
V_OTA_N_1903 PROBE<1903> VSS 0

* Device: OTA_P Size: 4 
V_OTA_P_1959 PROBE<1959> VSS 0
V_OTA_P_1960 PROBE<1960> VSS 0
V_OTA_P_1961 PROBE<1961> VDD 0
V_OTA_P_1962 PROBE<1962> VSS 0
V_OTA_P_1963 PROBE<1963> VSS 0

.ENDS

