
simulator lang=spice

.SUBCKT PK_NODE_external_connections 
+ NODE<1> NODE<2> NODE<3> NODE<4> NODE<5> 
+ NODE<6> NODE<7> NODE<8> NODE<9> NODE<10> 
+ NODE<11> NODE<12> NODE<13> NODE<14> NODE<15> 
+ NODE<16> NODE<17> NODE<18> NODE<19> NODE<20>        
+  pin<1> pin<2> pin<3> pin<4> pin<5> pin<6> pin<7>
+  pin<8> pin<9> pin<10> pin<11> pin<12> pin<13> pin<14> pin<15> pin<16> pin<17>
+  pin<18> pin<19> pin<20> pin<21> pin<22> pin<23> pin<24> pin<25> pin<26>
+  pin<27> pin<28> pin<29> pin<30> pin<31> pin<32> pin<33> pin<34> pin<35>
+  pin<36> pin<37> pin<38> pin<39> pin<40> pin<41> pin<42> pin<43> pin<44>
+  pin<45> pin<46> pin<47> pin<48> pin<49> pin<50> pin<51> pin<52> pin<53>
+  pin<54> pin<55> pin<56> pin<57> pin<58> pin<59> pin<60> pin<61> pin<62>
+  pin<63> pin<64> pin<65> pin<66> pin<67> pin<68> pin<69> pin<70> pin<71>
+  pin<72> pin<73> pin<74> pin<75> pin<76> pin<77> pin<78> pin<79> pin<80>
+  pin<81> pin<82> pin<83> pin<84> pin<85> pin<86> pin<87> pin<88> pin<89>
+  pin<90> pin<91> pin<92> pin<93> pin<94> pin<95> pin<96> pin<97> pin<98>
+  pin<99> pin<100>