
simulator lang=spice

.SUBCKT PK_set_sizes_2 PROBE<1889> PROBE<1890> PROBE<1891> PROBE<1892> PROBE<1893>
+  PROBE<1894> PROBE<1895> PROBE<1896> PROBE<1897> PROBE<1898> PROBE<1899>
+  PROBE<1900> PROBE<1901> PROBE<1902> PROBE<1903> PROBE<1904> PROBE<1905>
+  PROBE<1906> PROBE<1907> PROBE<1908> PROBE<1909> PROBE<1910> PROBE<1911>
+  PROBE<1912> PROBE<1913> PROBE<1914> PROBE<1915> PROBE<1916> PROBE<1917>
+  PROBE<1918> PROBE<1919> PROBE<1920> PROBE<1921> PROBE<1922> PROBE<1923>
+  PROBE<1924> PROBE<1925> PROBE<1926> PROBE<1927> PROBE<1928> PROBE<1929>
+  PROBE<1930> PROBE<1931> PROBE<1932> PROBE<1933> PROBE<1934> PROBE<1935>
+  PROBE<1936> PROBE<1937> PROBE<1938> PROBE<1939> PROBE<1940> PROBE<1941>
+  PROBE<1942> PROBE<1943> PROBE<1944> PROBE<1945> PROBE<1946> PROBE<1947>
+  PROBE<1948> PROBE<1949> PROBE<1950> PROBE<1951> PROBE<1952> PROBE<1953>
+  PROBE<1954> PROBE<1955> PROBE<1956> PROBE<1957> PROBE<1958> PROBE<1959>
+  PROBE<1960> PROBE<1961> PROBE<1962> PROBE<1963> PROBE<1964> PROBE<1965>
+  PROBE<1966> PROBE<1967> PROBE<1968> PROBE<1969> PROBE<1970> PROBE<1971>
+  PROBE<1972> PROBE<1973> PROBE<1974> PROBE<1975> PROBE<1976> PROBE<1977>
+  PROBE<1978> PROBE<1979> PROBE<1980> PROBE<1981> PROBE<1982> PROBE<1983>
+  PROBE<1984> PROBE<1985> PROBE<1986> PROBE<1987> PROBE<1988> PROBE<1989>
+  PROBE<1990> PROBE<1991> PROBE<1992> PROBE<1993> PROBE<1994> PROBE<1995>
+  PROBE<1996> PROBE<1997> PROBE<1998> PROBE<1999> PROBE<2000> PROBE<2001>
+  PROBE<2002> PROBE<2003> PROBE<2004> PROBE<2005> PROBE<2006> PROBE<2007>
+  PROBE<2008> VDD VSS